//	How to use:	
//	1. Edit the songs on the Enter Song sheet.	
// 	2. Select this whole worksheet, copy it, and paste it into a new file.	
//	3. Save the file as song_rom.v.	

module saw3_rom (
    input clk,						
	output reg [25:0] dout,						
	input [11:0] addr		
    );
        
    wire [25:0] memory [4095:0];  					
	always @(posedge clk)						
		dout = memory[addr];					

    parameter s1 = 142;
    parameter s2 = s1 + 646;
    parameter s3 = s2 + 81;

    assign memory[0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[79 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[80 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[81 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[82 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[83 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[84 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[85 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[86 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[87 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[88 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[89 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[90 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[91 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[92 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[93 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[94 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[95 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[96 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[97 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[98 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[99 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[100] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[101] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[102] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[103] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[104] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[105] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[106] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[107] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[108] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[109] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[110] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[111] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[112] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[113] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[114] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[115] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[116] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[117] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[118] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[119] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[120] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[121] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[122] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[123] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[124] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[125] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[126] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[127] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[128] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[129] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[130] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[131] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[132] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[133] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[134] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[135] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[136] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[137] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[138] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[139] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[140] = {7'd0  , 8'd123, 7'd0  , 2'd0, 2'd0};
    assign memory[141] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s1+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s1+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+25 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+26 ] = {7'd31 , 8'd96 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+27 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+28 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+29 ] = {7'd43 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+30 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+31 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+32 ] = {7'd31 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+33 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+34 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+35 ] = {7'd46 , 8'd96 , 7'd123, 2'd0, 2'd0};   //note: 5F#Gb
    assign memory[s1+36 ] = {7'd38 , 8'd96 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+37 ] = {7'd31 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+38 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+39 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+40 ] = {7'd43 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+41 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+42 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+43 ] = {7'd31 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+44 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+45 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+46 ] = {7'd46 , 8'd96 , 7'd123, 2'd0, 2'd0};   //note: 5F#Gb
    assign memory[s1+47 ] = {7'd38 , 8'd96 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+48 ] = {7'd31 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+49 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+50 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+51 ] = {7'd43 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+52 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+53 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+54 ] = {7'd31 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+55 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+56 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+57 ] = {7'd46 , 8'd96 , 7'd123, 2'd0, 2'd0};   //note: 5F#Gb
    assign memory[s1+58 ] = {7'd38 , 8'd96 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+59 ] = {7'd31 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+60 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+61 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+62 ] = {7'd43 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+63 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+64 ] = {7'd38 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+65 ] = {7'd31 , 8'd120, 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+67 ] = {7'd0  , 8'd9  , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+68 ] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+69 ] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+70 ] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+71 ] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+72 ] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+73 ] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+74 ] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+75 ] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+76 ] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+77 ] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+78 ] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+79 ] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+80 ] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+81 ] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+82 ] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+83 ] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+84 ] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+85 ] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+86 ] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+87 ] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+88 ] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+89 ] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+90 ] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+91 ] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+92 ] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+93 ] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+94 ] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+95 ] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+96 ] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+97 ] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+98 ] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+99 ] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+100] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+101] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+102] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+103] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+104] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+105] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+106] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+107] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+108] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+109] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+110] = {7'd30 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+111] = {7'd30 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+112] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+113] = {7'd42 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+114] = {7'd40 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+115] = {7'd42 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+116] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+117] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+118] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+119] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+120] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+121] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+122] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+123] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+124] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+125] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+126] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+127] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+128] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+129] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+130] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+131] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+132] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+133] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+134] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+135] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+136] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+137] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+138] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+139] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+140] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+141] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+142] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+143] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+144] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+145] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+146] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+147] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+148] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+149] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+150] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+151] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+152] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+153] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+154] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+155] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+156] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+157] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+158] = {7'd42 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+159] = {7'd42 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+160] = {7'd42 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+161] = {7'd42 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+162] = {7'd42 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+163] = {7'd42 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+164] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+165] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+166] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+167] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+168] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+169] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+170] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+171] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+172] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+173] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+174] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+175] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+176] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+177] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+178] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+179] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+180] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+181] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+182] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+183] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+184] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+185] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+186] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+187] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+188] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+189] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+190] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+191] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+192] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+193] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+194] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+195] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+196] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+197] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+198] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+199] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+200] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+201] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+202] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+203] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+204] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+205] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+206] = {7'd30 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+207] = {7'd30 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+208] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+209] = {7'd42 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+210] = {7'd40 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+211] = {7'd42 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+212] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+213] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+214] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+215] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+216] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+217] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+218] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+219] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+220] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+221] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+222] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+223] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+224] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+225] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+226] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+227] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+228] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+229] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+230] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+231] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+232] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+233] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+234] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+235] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+236] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+237] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+238] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+239] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+240] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+241] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+242] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+243] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+244] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+245] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+246] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+247] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+248] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+249] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+250] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+251] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+252] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+253] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+254] = {7'd30 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+255] = {7'd30 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+256] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+257] = {7'd42 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+258] = {7'd40 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+259] = {7'd42 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+260] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+261] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+262] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+263] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+264] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+265] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+266] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+267] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+268] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+269] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+270] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+271] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+272] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+273] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+274] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+275] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+276] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+277] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+278] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+279] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+280] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+281] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+282] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+283] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+284] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+285] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+286] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+287] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+288] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+289] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+290] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+291] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+292] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+293] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+294] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+295] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+296] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+297] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+298] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+299] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+300] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+301] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+302] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+303] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+304] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+305] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+306] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+307] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+308] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+309] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+310] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+311] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+312] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+313] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+314] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+315] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+316] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+317] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+318] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+319] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+320] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+321] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+322] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+323] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+324] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+325] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+326] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+327] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+328] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+329] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+330] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+331] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+332] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+333] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+334] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+335] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+336] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+337] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+338] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+339] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+340] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+341] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+342] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+343] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+344] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+345] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+346] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+347] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+348] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+349] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+350] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+351] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+352] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+353] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+354] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+355] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+356] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+357] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+358] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+359] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+360] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+361] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+362] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+363] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+364] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+365] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+366] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+367] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+368] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+369] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+370] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+371] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+372] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+373] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+374] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+375] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+376] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+377] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+378] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+379] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+380] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+381] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+382] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+383] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+384] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+385] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+386] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+387] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+388] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+389] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+390] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+391] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+392] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+393] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+394] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+395] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+396] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+397] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+398] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+399] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+400] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+401] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+402] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+403] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+404] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+405] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+406] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+407] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+408] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+409] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+410] = {7'd27 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+411] = {7'd27 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+412] = {7'd34 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+413] = {7'd39 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+414] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+415] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+416] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+417] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+418] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+419] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+420] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+421] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+422] = {7'd29 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+423] = {7'd29 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+424] = {7'd36 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+425] = {7'd41 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+426] = {7'd39 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+427] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+428] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+429] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+430] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+431] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+432] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+433] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+434] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+435] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+436] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+437] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+438] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+439] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+440] = {7'd31 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+441] = {7'd31 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+442] = {7'd38 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s1+443] = {7'd43 , 8'd48 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+444] = {7'd41 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+445] = {7'd43 , 8'd24 , 7'd113, 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+446] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+447] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+448] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+449] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+450] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+451] = {7'd31 , 8'd32 , 7'd113, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+452] = {7'd39 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s1+453] = {7'd39 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s1+454] = {7'd46 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5F#Gb
    assign memory[s1+455] = {7'd51 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+456] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+457] = {7'd51 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+458] = {7'd39 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s1+459] = {7'd39 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s1+460] = {7'd46 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5F#Gb
    assign memory[s1+461] = {7'd51 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+462] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+463] = {7'd51 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+464] = {7'd41 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+465] = {7'd41 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+466] = {7'd48 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5G#Ab
    assign memory[s1+467] = {7'd53 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+468] = {7'd51 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+469] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+470] = {7'd41 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+471] = {7'd41 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+472] = {7'd48 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5G#Ab
    assign memory[s1+473] = {7'd53 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+474] = {7'd51 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+475] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+476] = {7'd43 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+477] = {7'd43 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+478] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+479] = {7'd55 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+480] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+481] = {7'd55 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+482] = {7'd43 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+483] = {7'd43 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+484] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+485] = {7'd55 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+486] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+487] = {7'd55 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+488] = {7'd43 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+489] = {7'd43 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+490] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+491] = {7'd55 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+492] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+493] = {7'd55 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+494] = {7'd43 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+495] = {7'd43 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+496] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+497] = {7'd55 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+498] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+499] = {7'd55 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+500] = {7'd39 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s1+501] = {7'd39 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s1+502] = {7'd46 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5F#Gb
    assign memory[s1+503] = {7'd51 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+504] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+505] = {7'd51 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+506] = {7'd39 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s1+507] = {7'd39 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s1+508] = {7'd46 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5F#Gb
    assign memory[s1+509] = {7'd51 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+510] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+511] = {7'd51 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+512] = {7'd41 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+513] = {7'd41 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+514] = {7'd48 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5G#Ab
    assign memory[s1+515] = {7'd53 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+516] = {7'd51 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+517] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+518] = {7'd41 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+519] = {7'd41 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s1+520] = {7'd48 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5G#Ab
    assign memory[s1+521] = {7'd53 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+522] = {7'd51 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+523] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+524] = {7'd43 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+525] = {7'd43 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+526] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+527] = {7'd55 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+528] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+529] = {7'd55 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+530] = {7'd43 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+531] = {7'd43 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s1+532] = {7'd50 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 5A#Bb
    assign memory[s1+533] = {7'd55 , 8'd48 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+534] = {7'd53 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6C#Db
    assign memory[s1+535] = {7'd55 , 8'd24 , 7'd93 , 2'd0, 2'd0};   //note: 6D#Eb
    assign memory[s1+536] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+537] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+538] = {7'd28 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+539] = {7'd28 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+540] = {7'd35 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4G
    assign memory[s1+541] = {7'd40 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+542] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+543] = {7'd40 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+544] = {7'd28 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+545] = {7'd28 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+546] = {7'd35 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4G
    assign memory[s1+547] = {7'd40 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+548] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+549] = {7'd40 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+550] = {7'd30 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+551] = {7'd30 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+552] = {7'd37 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4A
    assign memory[s1+553] = {7'd42 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+554] = {7'd40 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+555] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+556] = {7'd30 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+557] = {7'd30 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+558] = {7'd37 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4A
    assign memory[s1+559] = {7'd42 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+560] = {7'd40 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+561] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+562] = {7'd32 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+563] = {7'd32 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+564] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+565] = {7'd44 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+566] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+567] = {7'd44 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+568] = {7'd32 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+569] = {7'd32 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+570] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+571] = {7'd44 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+572] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+573] = {7'd44 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+574] = {7'd32 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+575] = {7'd32 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+576] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+577] = {7'd44 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+578] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+579] = {7'd44 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+580] = {7'd32 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+581] = {7'd32 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+582] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+583] = {7'd44 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+584] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+585] = {7'd44 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+586] = {7'd28 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+587] = {7'd28 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+588] = {7'd35 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4G
    assign memory[s1+589] = {7'd40 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+590] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+591] = {7'd40 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+592] = {7'd28 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+593] = {7'd28 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+594] = {7'd35 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4G
    assign memory[s1+595] = {7'd40 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+596] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+597] = {7'd40 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+598] = {7'd30 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+599] = {7'd30 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+600] = {7'd37 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4A
    assign memory[s1+601] = {7'd42 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+602] = {7'd40 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+603] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+604] = {7'd30 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+605] = {7'd30 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+606] = {7'd37 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4A
    assign memory[s1+607] = {7'd42 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+608] = {7'd40 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5C
    assign memory[s1+609] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+610] = {7'd32 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+611] = {7'd32 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+612] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+613] = {7'd44 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+614] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+615] = {7'd44 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+616] = {7'd32 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+617] = {7'd32 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+618] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+619] = {7'd44 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+620] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+621] = {7'd44 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+622] = {7'd32 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+623] = {7'd32 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+624] = {7'd39 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4B
    assign memory[s1+625] = {7'd44 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+626] = {7'd42 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5D
    assign memory[s1+627] = {7'd44 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 5E
    assign memory[s1+628] = {7'd44 , 8'd48 , 7'd78 , 2'd0, 2'd0};   //note: 5E
    assign memory[s1+629] = {7'd44 , 8'd24 , 7'd78 , 2'd0, 2'd0};   //note: 5E
    assign memory[s1+630] = {7'd51 , 8'd24 , 7'd78 , 2'd0, 2'd0};   //note: 5B
    assign memory[s1+631] = {7'd56 , 8'd48 , 7'd78 , 2'd0, 2'd0};   //note: 6E
    assign memory[s1+632] = {7'd54 , 8'd24 , 7'd78 , 2'd0, 2'd0};   //note: 6D
    assign memory[s1+633] = {7'd56 , 8'd24 , 7'd78 , 2'd0, 2'd0};   //note: 6E
    assign memory[s1+634] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+635] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+636] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+637] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+638] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+639] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+640] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+641] = {7'd0  , 8'd135, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+642] = {7'd0  , 8'd1  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+643] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+644] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+645] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s2+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s2+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+79 ] = {7'd0  , 8'd79 , 7'd0  , 2'd0, 2'd0};
    assign memory[s2+80 ] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s3+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s3+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+74 ] = {7'd0  , 8'd107, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+75 ] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

endmodule							
