`timescale 1ns / 1ps
module number_rom_reader(
    input clk,
    input [9:0]progress,
    input [4:0]x1,
    input [4:0]x2,
    input [4:0]x3,
    input [4:0]y,
    output [1:0] ui_pixel_type1,
    output [1:0] ui_pixel_type2,
    output [1:0] ui_pixel_type3
    );

    wire [3:0] prog1, prog2, prog3;
    wire [1:0] ui_pixel_type1_mid;
    assign ui_pixel_type1 = ui_pixel_type1_mid & {1'd0,prog1!=0};
    assign prog3 = progress % 10;
    assign prog2 = progress / 10 % 10;
    assign prog1 = (progress>=1000) ? 0 : progress / 100;

    wire [12:0] nbr_in1,nbr_in2,nbr_in3;

    assign nbr_in1 = 180*y+18*prog1+x1;
    assign nbr_in2 = 180*y+18*prog2+x2;
    assign nbr_in3 = 180*y+18*prog3+x3;
    number_rom nbr1(
        .clk        (clk),
        .nbr_in      (nbr_in1),
        .dout       (ui_pixel_type1_mid)
    );
    number_rom nbr2(
        .clk        (clk)   , 
        .nbr_in      (nbr_in2),
        .dout       (ui_pixel_type2)
    );
    number_rom nbr3(
        .clk        (clk),    
        .nbr_in      (nbr_in3),
        .dout       (ui_pixel_type3)
    );

endmodule
module number_rom(
    input clk,
    input [12:0]nbr_in,
    output reg[1:0] dout
    );
    wire [1:0] memnumber [4319:0];
    always @(posedge clk)begin
        dout = memnumber [nbr_in];
    end
    
    
    
    assign memnumber[0   ] = 2'd0;
    assign memnumber[1   ] = 2'd0;
    assign memnumber[2   ] = 2'd0;
    assign memnumber[3   ] = 2'd0;
    assign memnumber[4   ] = 2'd0;
    assign memnumber[5   ] = 2'd2;
    assign memnumber[6   ] = 2'd2;
    assign memnumber[7   ] = 2'd2;
    assign memnumber[8   ] = 2'd2;
    assign memnumber[9   ] = 2'd2;
    assign memnumber[10  ] = 2'd2;
    assign memnumber[11  ] = 2'd0;
    assign memnumber[12  ] = 2'd0;
    assign memnumber[13  ] = 2'd0;
    assign memnumber[14  ] = 2'd0;
    assign memnumber[15  ] = 2'd0;
    assign memnumber[16  ] = 2'd0;
    assign memnumber[17  ] = 2'd0;
    assign memnumber[18  ] = 2'd0;
    assign memnumber[19  ] = 2'd0;
    assign memnumber[20  ] = 2'd0;
    assign memnumber[21  ] = 2'd0;
    assign memnumber[22  ] = 2'd0;
    assign memnumber[23  ] = 2'd2;
    assign memnumber[24  ] = 2'd2;
    assign memnumber[25  ] = 2'd2;
    assign memnumber[26  ] = 2'd2;
    assign memnumber[27  ] = 2'd2;
    assign memnumber[28  ] = 2'd0;
    assign memnumber[29  ] = 2'd0;
    assign memnumber[30  ] = 2'd0;
    assign memnumber[31  ] = 2'd0;
    assign memnumber[32  ] = 2'd0;
    assign memnumber[33  ] = 2'd0;
    assign memnumber[34  ] = 2'd0;
    assign memnumber[35  ] = 2'd0;
    assign memnumber[36  ] = 2'd0;
    assign memnumber[37  ] = 2'd0;
    assign memnumber[38  ] = 2'd0;
    assign memnumber[39  ] = 2'd0;
    assign memnumber[40  ] = 2'd0;
    assign memnumber[41  ] = 2'd0;
    assign memnumber[42  ] = 2'd2;
    assign memnumber[43  ] = 2'd2;
    assign memnumber[44  ] = 2'd2;
    assign memnumber[45  ] = 2'd2;
    assign memnumber[46  ] = 2'd2;
    assign memnumber[47  ] = 2'd2;
    assign memnumber[48  ] = 2'd0;
    assign memnumber[49  ] = 2'd0;
    assign memnumber[50  ] = 2'd0;
    assign memnumber[51  ] = 2'd0;
    assign memnumber[52  ] = 2'd0;
    assign memnumber[53  ] = 2'd0;
    assign memnumber[54  ] = 2'd0;
    assign memnumber[55  ] = 2'd0;
    assign memnumber[56  ] = 2'd0;
    assign memnumber[57  ] = 2'd0;
    assign memnumber[58  ] = 2'd0;
    assign memnumber[59  ] = 2'd2;
    assign memnumber[60  ] = 2'd2;
    assign memnumber[61  ] = 2'd2;
    assign memnumber[62  ] = 2'd2;
    assign memnumber[63  ] = 2'd2;
    assign memnumber[64  ] = 2'd2;
    assign memnumber[65  ] = 2'd0;
    assign memnumber[66  ] = 2'd0;
    assign memnumber[67  ] = 2'd0;
    assign memnumber[68  ] = 2'd0;
    assign memnumber[69  ] = 2'd0;
    assign memnumber[70  ] = 2'd0;
    assign memnumber[71  ] = 2'd0;
    assign memnumber[72  ] = 2'd0;
    assign memnumber[73  ] = 2'd0;
    assign memnumber[74  ] = 2'd0;
    assign memnumber[75  ] = 2'd0;
    assign memnumber[76  ] = 2'd0;
    assign memnumber[77  ] = 2'd0;
    assign memnumber[78  ] = 2'd0;
    assign memnumber[79  ] = 2'd0;
    assign memnumber[80  ] = 2'd0;
    assign memnumber[81  ] = 2'd0;
    assign memnumber[82  ] = 2'd0;
    assign memnumber[83  ] = 2'd0;
    assign memnumber[84  ] = 2'd2;
    assign memnumber[85  ] = 2'd0;
    assign memnumber[86  ] = 2'd0;
    assign memnumber[87  ] = 2'd0;
    assign memnumber[88  ] = 2'd0;
    assign memnumber[89  ] = 2'd0;
    assign memnumber[90  ] = 2'd0;
    assign memnumber[91  ] = 2'd0;
    assign memnumber[92  ] = 2'd0;
    assign memnumber[93  ] = 2'd0;
    assign memnumber[94  ] = 2'd2;
    assign memnumber[95  ] = 2'd2;
    assign memnumber[96  ] = 2'd2;
    assign memnumber[97  ] = 2'd2;
    assign memnumber[98  ] = 2'd2;
    assign memnumber[99  ] = 2'd2;
    assign memnumber[100 ] = 2'd2;
    assign memnumber[101 ] = 2'd2;
    assign memnumber[102 ] = 2'd2;
    assign memnumber[103 ] = 2'd2;
    assign memnumber[104 ] = 2'd0;
    assign memnumber[105 ] = 2'd0;
    assign memnumber[106 ] = 2'd0;
    assign memnumber[107 ] = 2'd0;
    assign memnumber[108 ] = 2'd0;
    assign memnumber[109 ] = 2'd0;
    assign memnumber[110 ] = 2'd0;
    assign memnumber[111 ] = 2'd0;
    assign memnumber[112 ] = 2'd0;
    assign memnumber[113 ] = 2'd0;
    assign memnumber[114 ] = 2'd0;
    assign memnumber[115 ] = 2'd0;
    assign memnumber[116 ] = 2'd0;
    assign memnumber[117 ] = 2'd0;
    assign memnumber[118 ] = 2'd2;
    assign memnumber[119 ] = 2'd2;
    assign memnumber[120 ] = 2'd0;
    assign memnumber[121 ] = 2'd0;
    assign memnumber[122 ] = 2'd0;
    assign memnumber[123 ] = 2'd0;
    assign memnumber[124 ] = 2'd0;
    assign memnumber[125 ] = 2'd0;
    assign memnumber[126 ] = 2'd0;
    assign memnumber[127 ] = 2'd0;
    assign memnumber[128 ] = 2'd2;
    assign memnumber[129 ] = 2'd2;
    assign memnumber[130 ] = 2'd2;
    assign memnumber[131 ] = 2'd2;
    assign memnumber[132 ] = 2'd2;
    assign memnumber[133 ] = 2'd2;
    assign memnumber[134 ] = 2'd2;
    assign memnumber[135 ] = 2'd2;
    assign memnumber[136 ] = 2'd2;
    assign memnumber[137 ] = 2'd2;
    assign memnumber[138 ] = 2'd2;
    assign memnumber[139 ] = 2'd2;
    assign memnumber[140 ] = 2'd2;
    assign memnumber[141 ] = 2'd2;
    assign memnumber[142 ] = 2'd0;
    assign memnumber[143 ] = 2'd0;
    assign memnumber[144 ] = 2'd0;
    assign memnumber[145 ] = 2'd0;
    assign memnumber[146 ] = 2'd0;
    assign memnumber[147 ] = 2'd0;
    assign memnumber[148 ] = 2'd0;
    assign memnumber[149 ] = 2'd2;
    assign memnumber[150 ] = 2'd2;
    assign memnumber[151 ] = 2'd2;
    assign memnumber[152 ] = 2'd2;
    assign memnumber[153 ] = 2'd2;
    assign memnumber[154 ] = 2'd2;
    assign memnumber[155 ] = 2'd0;
    assign memnumber[156 ] = 2'd0;
    assign memnumber[157 ] = 2'd0;
    assign memnumber[158 ] = 2'd0;
    assign memnumber[159 ] = 2'd0;
    assign memnumber[160 ] = 2'd0;
    assign memnumber[161 ] = 2'd0;
    assign memnumber[162 ] = 2'd0;
    assign memnumber[163 ] = 2'd0;
    assign memnumber[164 ] = 2'd0;
    assign memnumber[165 ] = 2'd0;
    assign memnumber[166 ] = 2'd0;
    assign memnumber[167 ] = 2'd2;
    assign memnumber[168 ] = 2'd2;
    assign memnumber[169 ] = 2'd2;
    assign memnumber[170 ] = 2'd2;
    assign memnumber[171 ] = 2'd2;
    assign memnumber[172 ] = 2'd0;
    assign memnumber[173 ] = 2'd0;
    assign memnumber[174 ] = 2'd0;
    assign memnumber[175 ] = 2'd0;
    assign memnumber[176 ] = 2'd0;
    assign memnumber[177 ] = 2'd0;
    assign memnumber[178 ] = 2'd0;
    assign memnumber[179 ] = 2'd0;
    assign memnumber[180 ] = 2'd0;
    assign memnumber[181 ] = 2'd0;
    assign memnumber[182 ] = 2'd0;
    assign memnumber[183 ] = 2'd2;
    assign memnumber[184 ] = 2'd2;
    assign memnumber[185 ] = 2'd2;
    assign memnumber[186 ] = 2'd2;
    assign memnumber[187 ] = 2'd2;
    assign memnumber[188 ] = 2'd2;
    assign memnumber[189 ] = 2'd2;
    assign memnumber[190 ] = 2'd2;
    assign memnumber[191 ] = 2'd2;
    assign memnumber[192 ] = 2'd0;
    assign memnumber[193 ] = 2'd0;
    assign memnumber[194 ] = 2'd0;
    assign memnumber[195 ] = 2'd0;
    assign memnumber[196 ] = 2'd0;
    assign memnumber[197 ] = 2'd0;
    assign memnumber[198 ] = 2'd0;
    assign memnumber[199 ] = 2'd0;
    assign memnumber[200 ] = 2'd0;
    assign memnumber[201 ] = 2'd0;
    assign memnumber[202 ] = 2'd2;
    assign memnumber[203 ] = 2'd2;
    assign memnumber[204 ] = 2'd2;
    assign memnumber[205 ] = 2'd2;
    assign memnumber[206 ] = 2'd2;
    assign memnumber[207 ] = 2'd2;
    assign memnumber[208 ] = 2'd1;
    assign memnumber[209 ] = 2'd0;
    assign memnumber[210 ] = 2'd0;
    assign memnumber[211 ] = 2'd0;
    assign memnumber[212 ] = 2'd0;
    assign memnumber[213 ] = 2'd0;
    assign memnumber[214 ] = 2'd0;
    assign memnumber[215 ] = 2'd0;
    assign memnumber[216 ] = 2'd0;
    assign memnumber[217 ] = 2'd0;
    assign memnumber[218 ] = 2'd0;
    assign memnumber[219 ] = 2'd0;
    assign memnumber[220 ] = 2'd2;
    assign memnumber[221 ] = 2'd2;
    assign memnumber[222 ] = 2'd2;
    assign memnumber[223 ] = 2'd2;
    assign memnumber[224 ] = 2'd2;
    assign memnumber[225 ] = 2'd2;
    assign memnumber[226 ] = 2'd2;
    assign memnumber[227 ] = 2'd2;
    assign memnumber[228 ] = 2'd2;
    assign memnumber[229 ] = 2'd0;
    assign memnumber[230 ] = 2'd0;
    assign memnumber[231 ] = 2'd0;
    assign memnumber[232 ] = 2'd0;
    assign memnumber[233 ] = 2'd0;
    assign memnumber[234 ] = 2'd0;
    assign memnumber[235 ] = 2'd0;
    assign memnumber[236 ] = 2'd0;
    assign memnumber[237 ] = 2'd0;
    assign memnumber[238 ] = 2'd2;
    assign memnumber[239 ] = 2'd2;
    assign memnumber[240 ] = 2'd2;
    assign memnumber[241 ] = 2'd2;
    assign memnumber[242 ] = 2'd2;
    assign memnumber[243 ] = 2'd2;
    assign memnumber[244 ] = 2'd2;
    assign memnumber[245 ] = 2'd2;
    assign memnumber[246 ] = 2'd2;
    assign memnumber[247 ] = 2'd0;
    assign memnumber[248 ] = 2'd0;
    assign memnumber[249 ] = 2'd0;
    assign memnumber[250 ] = 2'd0;
    assign memnumber[251 ] = 2'd0;
    assign memnumber[252 ] = 2'd0;
    assign memnumber[253 ] = 2'd0;
    assign memnumber[254 ] = 2'd0;
    assign memnumber[255 ] = 2'd0;
    assign memnumber[256 ] = 2'd0;
    assign memnumber[257 ] = 2'd0;
    assign memnumber[258 ] = 2'd0;
    assign memnumber[259 ] = 2'd0;
    assign memnumber[260 ] = 2'd0;
    assign memnumber[261 ] = 2'd0;
    assign memnumber[262 ] = 2'd0;
    assign memnumber[263 ] = 2'd0;
    assign memnumber[264 ] = 2'd2;
    assign memnumber[265 ] = 2'd1;
    assign memnumber[266 ] = 2'd0;
    assign memnumber[267 ] = 2'd0;
    assign memnumber[268 ] = 2'd0;
    assign memnumber[269 ] = 2'd0;
    assign memnumber[270 ] = 2'd0;
    assign memnumber[271 ] = 2'd0;
    assign memnumber[272 ] = 2'd0;
    assign memnumber[273 ] = 2'd0;
    assign memnumber[274 ] = 2'd2;
    assign memnumber[275 ] = 2'd2;
    assign memnumber[276 ] = 2'd2;
    assign memnumber[277 ] = 2'd2;
    assign memnumber[278 ] = 2'd2;
    assign memnumber[279 ] = 2'd2;
    assign memnumber[280 ] = 2'd2;
    assign memnumber[281 ] = 2'd2;
    assign memnumber[282 ] = 2'd2;
    assign memnumber[283 ] = 2'd2;
    assign memnumber[284 ] = 2'd1;
    assign memnumber[285 ] = 2'd0;
    assign memnumber[286 ] = 2'd0;
    assign memnumber[287 ] = 2'd0;
    assign memnumber[288 ] = 2'd0;
    assign memnumber[289 ] = 2'd0;
    assign memnumber[290 ] = 2'd0;
    assign memnumber[291 ] = 2'd0;
    assign memnumber[292 ] = 2'd0;
    assign memnumber[293 ] = 2'd0;
    assign memnumber[294 ] = 2'd0;
    assign memnumber[295 ] = 2'd0;
    assign memnumber[296 ] = 2'd0;
    assign memnumber[297 ] = 2'd2;
    assign memnumber[298 ] = 2'd2;
    assign memnumber[299 ] = 2'd1;
    assign memnumber[300 ] = 2'd1;
    assign memnumber[301 ] = 2'd0;
    assign memnumber[302 ] = 2'd0;
    assign memnumber[303 ] = 2'd0;
    assign memnumber[304 ] = 2'd0;
    assign memnumber[305 ] = 2'd0;
    assign memnumber[306 ] = 2'd0;
    assign memnumber[307 ] = 2'd0;
    assign memnumber[308 ] = 2'd2;
    assign memnumber[309 ] = 2'd2;
    assign memnumber[310 ] = 2'd2;
    assign memnumber[311 ] = 2'd2;
    assign memnumber[312 ] = 2'd2;
    assign memnumber[313 ] = 2'd2;
    assign memnumber[314 ] = 2'd2;
    assign memnumber[315 ] = 2'd2;
    assign memnumber[316 ] = 2'd2;
    assign memnumber[317 ] = 2'd2;
    assign memnumber[318 ] = 2'd2;
    assign memnumber[319 ] = 2'd2;
    assign memnumber[320 ] = 2'd2;
    assign memnumber[321 ] = 2'd1;
    assign memnumber[322 ] = 2'd1;
    assign memnumber[323 ] = 2'd0;
    assign memnumber[324 ] = 2'd0;
    assign memnumber[325 ] = 2'd0;
    assign memnumber[326 ] = 2'd0;
    assign memnumber[327 ] = 2'd2;
    assign memnumber[328 ] = 2'd2;
    assign memnumber[329 ] = 2'd2;
    assign memnumber[330 ] = 2'd2;
    assign memnumber[331 ] = 2'd2;
    assign memnumber[332 ] = 2'd2;
    assign memnumber[333 ] = 2'd2;
    assign memnumber[334 ] = 2'd2;
    assign memnumber[335 ] = 2'd2;
    assign memnumber[336 ] = 2'd2;
    assign memnumber[337 ] = 2'd0;
    assign memnumber[338 ] = 2'd0;
    assign memnumber[339 ] = 2'd0;
    assign memnumber[340 ] = 2'd0;
    assign memnumber[341 ] = 2'd0;
    assign memnumber[342 ] = 2'd0;
    assign memnumber[343 ] = 2'd0;
    assign memnumber[344 ] = 2'd0;
    assign memnumber[345 ] = 2'd2;
    assign memnumber[346 ] = 2'd2;
    assign memnumber[347 ] = 2'd2;
    assign memnumber[348 ] = 2'd2;
    assign memnumber[349 ] = 2'd2;
    assign memnumber[350 ] = 2'd2;
    assign memnumber[351 ] = 2'd2;
    assign memnumber[352 ] = 2'd2;
    assign memnumber[353 ] = 2'd2;
    assign memnumber[354 ] = 2'd0;
    assign memnumber[355 ] = 2'd0;
    assign memnumber[356 ] = 2'd0;
    assign memnumber[357 ] = 2'd0;
    assign memnumber[358 ] = 2'd0;
    assign memnumber[359 ] = 2'd0;
    assign memnumber[360 ] = 2'd0;
    assign memnumber[361 ] = 2'd0;
    assign memnumber[362 ] = 2'd2;
    assign memnumber[363 ] = 2'd2;
    assign memnumber[364 ] = 2'd2;
    assign memnumber[365 ] = 2'd2;
    assign memnumber[366 ] = 2'd1;
    assign memnumber[367 ] = 2'd1;
    assign memnumber[368 ] = 2'd1;
    assign memnumber[369 ] = 2'd1;
    assign memnumber[370 ] = 2'd2;
    assign memnumber[371 ] = 2'd2;
    assign memnumber[372 ] = 2'd2;
    assign memnumber[373 ] = 2'd0;
    assign memnumber[374 ] = 2'd0;
    assign memnumber[375 ] = 2'd0;
    assign memnumber[376 ] = 2'd0;
    assign memnumber[377 ] = 2'd0;
    assign memnumber[378 ] = 2'd0;
    assign memnumber[379 ] = 2'd0;
    assign memnumber[380 ] = 2'd0;
    assign memnumber[381 ] = 2'd0;
    assign memnumber[382 ] = 2'd0;
    assign memnumber[383 ] = 2'd1;
    assign memnumber[384 ] = 2'd1;
    assign memnumber[385 ] = 2'd1;
    assign memnumber[386 ] = 2'd2;
    assign memnumber[387 ] = 2'd2;
    assign memnumber[388 ] = 2'd1;
    assign memnumber[389 ] = 2'd0;
    assign memnumber[390 ] = 2'd0;
    assign memnumber[391 ] = 2'd0;
    assign memnumber[392 ] = 2'd0;
    assign memnumber[393 ] = 2'd0;
    assign memnumber[394 ] = 2'd0;
    assign memnumber[395 ] = 2'd0;
    assign memnumber[396 ] = 2'd0;
    assign memnumber[397 ] = 2'd0;
    assign memnumber[398 ] = 2'd0;
    assign memnumber[399 ] = 2'd2;
    assign memnumber[400 ] = 2'd2;
    assign memnumber[401 ] = 2'd2;
    assign memnumber[402 ] = 2'd1;
    assign memnumber[403 ] = 2'd1;
    assign memnumber[404 ] = 2'd1;
    assign memnumber[405 ] = 2'd1;
    assign memnumber[406 ] = 2'd1;
    assign memnumber[407 ] = 2'd2;
    assign memnumber[408 ] = 2'd2;
    assign memnumber[409 ] = 2'd2;
    assign memnumber[410 ] = 2'd0;
    assign memnumber[411 ] = 2'd0;
    assign memnumber[412 ] = 2'd0;
    assign memnumber[413 ] = 2'd0;
    assign memnumber[414 ] = 2'd0;
    assign memnumber[415 ] = 2'd0;
    assign memnumber[416 ] = 2'd0;
    assign memnumber[417 ] = 2'd2;
    assign memnumber[418 ] = 2'd2;
    assign memnumber[419 ] = 2'd2;
    assign memnumber[420 ] = 2'd1;
    assign memnumber[421 ] = 2'd1;
    assign memnumber[422 ] = 2'd1;
    assign memnumber[423 ] = 2'd1;
    assign memnumber[424 ] = 2'd1;
    assign memnumber[425 ] = 2'd2;
    assign memnumber[426 ] = 2'd2;
    assign memnumber[427 ] = 2'd2;
    assign memnumber[428 ] = 2'd0;
    assign memnumber[429 ] = 2'd0;
    assign memnumber[430 ] = 2'd0;
    assign memnumber[431 ] = 2'd0;
    assign memnumber[432 ] = 2'd0;
    assign memnumber[433 ] = 2'd0;
    assign memnumber[434 ] = 2'd0;
    assign memnumber[435 ] = 2'd0;
    assign memnumber[436 ] = 2'd0;
    assign memnumber[437 ] = 2'd0;
    assign memnumber[438 ] = 2'd0;
    assign memnumber[439 ] = 2'd0;
    assign memnumber[440 ] = 2'd0;
    assign memnumber[441 ] = 2'd0;
    assign memnumber[442 ] = 2'd0;
    assign memnumber[443 ] = 2'd2;
    assign memnumber[444 ] = 2'd2;
    assign memnumber[445 ] = 2'd1;
    assign memnumber[446 ] = 2'd0;
    assign memnumber[447 ] = 2'd0;
    assign memnumber[448 ] = 2'd0;
    assign memnumber[449 ] = 2'd0;
    assign memnumber[450 ] = 2'd0;
    assign memnumber[451 ] = 2'd0;
    assign memnumber[452 ] = 2'd0;
    assign memnumber[453 ] = 2'd0;
    assign memnumber[454 ] = 2'd2;
    assign memnumber[455 ] = 2'd2;
    assign memnumber[456 ] = 2'd1;
    assign memnumber[457 ] = 2'd1;
    assign memnumber[458 ] = 2'd1;
    assign memnumber[459 ] = 2'd1;
    assign memnumber[460 ] = 2'd1;
    assign memnumber[461 ] = 2'd1;
    assign memnumber[462 ] = 2'd1;
    assign memnumber[463 ] = 2'd1;
    assign memnumber[464 ] = 2'd1;
    assign memnumber[465 ] = 2'd0;
    assign memnumber[466 ] = 2'd0;
    assign memnumber[467 ] = 2'd0;
    assign memnumber[468 ] = 2'd0;
    assign memnumber[469 ] = 2'd0;
    assign memnumber[470 ] = 2'd0;
    assign memnumber[471 ] = 2'd0;
    assign memnumber[472 ] = 2'd0;
    assign memnumber[473 ] = 2'd0;
    assign memnumber[474 ] = 2'd0;
    assign memnumber[475 ] = 2'd0;
    assign memnumber[476 ] = 2'd2;
    assign memnumber[477 ] = 2'd2;
    assign memnumber[478 ] = 2'd2;
    assign memnumber[479 ] = 2'd1;
    assign memnumber[480 ] = 2'd0;
    assign memnumber[481 ] = 2'd0;
    assign memnumber[482 ] = 2'd0;
    assign memnumber[483 ] = 2'd0;
    assign memnumber[484 ] = 2'd0;
    assign memnumber[485 ] = 2'd0;
    assign memnumber[486 ] = 2'd0;
    assign memnumber[487 ] = 2'd0;
    assign memnumber[488 ] = 2'd0;
    assign memnumber[489 ] = 2'd1;
    assign memnumber[490 ] = 2'd1;
    assign memnumber[491 ] = 2'd1;
    assign memnumber[492 ] = 2'd1;
    assign memnumber[493 ] = 2'd1;
    assign memnumber[494 ] = 2'd1;
    assign memnumber[495 ] = 2'd1;
    assign memnumber[496 ] = 2'd1;
    assign memnumber[497 ] = 2'd1;
    assign memnumber[498 ] = 2'd1;
    assign memnumber[499 ] = 2'd2;
    assign memnumber[500 ] = 2'd2;
    assign memnumber[501 ] = 2'd1;
    assign memnumber[502 ] = 2'd0;
    assign memnumber[503 ] = 2'd0;
    assign memnumber[504 ] = 2'd0;
    assign memnumber[505 ] = 2'd0;
    assign memnumber[506 ] = 2'd2;
    assign memnumber[507 ] = 2'd2;
    assign memnumber[508 ] = 2'd2;
    assign memnumber[509 ] = 2'd1;
    assign memnumber[510 ] = 2'd1;
    assign memnumber[511 ] = 2'd1;
    assign memnumber[512 ] = 2'd1;
    assign memnumber[513 ] = 2'd1;
    assign memnumber[514 ] = 2'd1;
    assign memnumber[515 ] = 2'd2;
    assign memnumber[516 ] = 2'd2;
    assign memnumber[517 ] = 2'd2;
    assign memnumber[518 ] = 2'd0;
    assign memnumber[519 ] = 2'd0;
    assign memnumber[520 ] = 2'd0;
    assign memnumber[521 ] = 2'd0;
    assign memnumber[522 ] = 2'd0;
    assign memnumber[523 ] = 2'd0;
    assign memnumber[524 ] = 2'd2;
    assign memnumber[525 ] = 2'd2;
    assign memnumber[526 ] = 2'd2;
    assign memnumber[527 ] = 2'd1;
    assign memnumber[528 ] = 2'd1;
    assign memnumber[529 ] = 2'd1;
    assign memnumber[530 ] = 2'd1;
    assign memnumber[531 ] = 2'd1;
    assign memnumber[532 ] = 2'd2;
    assign memnumber[533 ] = 2'd2;
    assign memnumber[534 ] = 2'd2;
    assign memnumber[535 ] = 2'd0;
    assign memnumber[536 ] = 2'd0;
    assign memnumber[537 ] = 2'd0;
    assign memnumber[538 ] = 2'd0;
    assign memnumber[539 ] = 2'd0;
    assign memnumber[540 ] = 2'd0;
    assign memnumber[541 ] = 2'd0;
    assign memnumber[542 ] = 2'd2;
    assign memnumber[543 ] = 2'd2;
    assign memnumber[544 ] = 2'd1;
    assign memnumber[545 ] = 2'd1;
    assign memnumber[546 ] = 2'd1;
    assign memnumber[547 ] = 2'd0;
    assign memnumber[548 ] = 2'd0;
    assign memnumber[549 ] = 2'd0;
    assign memnumber[550 ] = 2'd0;
    assign memnumber[551 ] = 2'd1;
    assign memnumber[552 ] = 2'd2;
    assign memnumber[553 ] = 2'd2;
    assign memnumber[554 ] = 2'd0;
    assign memnumber[555 ] = 2'd0;
    assign memnumber[556 ] = 2'd0;
    assign memnumber[557 ] = 2'd0;
    assign memnumber[558 ] = 2'd0;
    assign memnumber[559 ] = 2'd0;
    assign memnumber[560 ] = 2'd0;
    assign memnumber[561 ] = 2'd0;
    assign memnumber[562 ] = 2'd0;
    assign memnumber[563 ] = 2'd0;
    assign memnumber[564 ] = 2'd0;
    assign memnumber[565 ] = 2'd0;
    assign memnumber[566 ] = 2'd2;
    assign memnumber[567 ] = 2'd2;
    assign memnumber[568 ] = 2'd1;
    assign memnumber[569 ] = 2'd0;
    assign memnumber[570 ] = 2'd0;
    assign memnumber[571 ] = 2'd0;
    assign memnumber[572 ] = 2'd0;
    assign memnumber[573 ] = 2'd0;
    assign memnumber[574 ] = 2'd0;
    assign memnumber[575 ] = 2'd0;
    assign memnumber[576 ] = 2'd0;
    assign memnumber[577 ] = 2'd0;
    assign memnumber[578 ] = 2'd2;
    assign memnumber[579 ] = 2'd2;
    assign memnumber[580 ] = 2'd2;
    assign memnumber[581 ] = 2'd1;
    assign memnumber[582 ] = 2'd1;
    assign memnumber[583 ] = 2'd0;
    assign memnumber[584 ] = 2'd0;
    assign memnumber[585 ] = 2'd0;
    assign memnumber[586 ] = 2'd0;
    assign memnumber[587 ] = 2'd0;
    assign memnumber[588 ] = 2'd1;
    assign memnumber[589 ] = 2'd2;
    assign memnumber[590 ] = 2'd2;
    assign memnumber[591 ] = 2'd0;
    assign memnumber[592 ] = 2'd0;
    assign memnumber[593 ] = 2'd0;
    assign memnumber[594 ] = 2'd0;
    assign memnumber[595 ] = 2'd0;
    assign memnumber[596 ] = 2'd2;
    assign memnumber[597 ] = 2'd2;
    assign memnumber[598 ] = 2'd1;
    assign memnumber[599 ] = 2'd1;
    assign memnumber[600 ] = 2'd1;
    assign memnumber[601 ] = 2'd0;
    assign memnumber[602 ] = 2'd0;
    assign memnumber[603 ] = 2'd0;
    assign memnumber[604 ] = 2'd0;
    assign memnumber[605 ] = 2'd0;
    assign memnumber[606 ] = 2'd2;
    assign memnumber[607 ] = 2'd2;
    assign memnumber[608 ] = 2'd2;
    assign memnumber[609 ] = 2'd0;
    assign memnumber[610 ] = 2'd0;
    assign memnumber[611 ] = 2'd0;
    assign memnumber[612 ] = 2'd0;
    assign memnumber[613 ] = 2'd0;
    assign memnumber[614 ] = 2'd0;
    assign memnumber[615 ] = 2'd0;
    assign memnumber[616 ] = 2'd0;
    assign memnumber[617 ] = 2'd0;
    assign memnumber[618 ] = 2'd0;
    assign memnumber[619 ] = 2'd0;
    assign memnumber[620 ] = 2'd0;
    assign memnumber[621 ] = 2'd0;
    assign memnumber[622 ] = 2'd2;
    assign memnumber[623 ] = 2'd2;
    assign memnumber[624 ] = 2'd2;
    assign memnumber[625 ] = 2'd1;
    assign memnumber[626 ] = 2'd0;
    assign memnumber[627 ] = 2'd0;
    assign memnumber[628 ] = 2'd0;
    assign memnumber[629 ] = 2'd0;
    assign memnumber[630 ] = 2'd0;
    assign memnumber[631 ] = 2'd0;
    assign memnumber[632 ] = 2'd0;
    assign memnumber[633 ] = 2'd2;
    assign memnumber[634 ] = 2'd2;
    assign memnumber[635 ] = 2'd1;
    assign memnumber[636 ] = 2'd1;
    assign memnumber[637 ] = 2'd0;
    assign memnumber[638 ] = 2'd0;
    assign memnumber[639 ] = 2'd0;
    assign memnumber[640 ] = 2'd0;
    assign memnumber[641 ] = 2'd0;
    assign memnumber[642 ] = 2'd0;
    assign memnumber[643 ] = 2'd0;
    assign memnumber[644 ] = 2'd0;
    assign memnumber[645 ] = 2'd0;
    assign memnumber[646 ] = 2'd0;
    assign memnumber[647 ] = 2'd0;
    assign memnumber[648 ] = 2'd0;
    assign memnumber[649 ] = 2'd0;
    assign memnumber[650 ] = 2'd0;
    assign memnumber[651 ] = 2'd0;
    assign memnumber[652 ] = 2'd0;
    assign memnumber[653 ] = 2'd0;
    assign memnumber[654 ] = 2'd0;
    assign memnumber[655 ] = 2'd0;
    assign memnumber[656 ] = 2'd2;
    assign memnumber[657 ] = 2'd2;
    assign memnumber[658 ] = 2'd1;
    assign memnumber[659 ] = 2'd1;
    assign memnumber[660 ] = 2'd0;
    assign memnumber[661 ] = 2'd0;
    assign memnumber[662 ] = 2'd0;
    assign memnumber[663 ] = 2'd0;
    assign memnumber[664 ] = 2'd0;
    assign memnumber[665 ] = 2'd0;
    assign memnumber[666 ] = 2'd0;
    assign memnumber[667 ] = 2'd0;
    assign memnumber[668 ] = 2'd0;
    assign memnumber[669 ] = 2'd0;
    assign memnumber[670 ] = 2'd0;
    assign memnumber[671 ] = 2'd0;
    assign memnumber[672 ] = 2'd0;
    assign memnumber[673 ] = 2'd0;
    assign memnumber[674 ] = 2'd0;
    assign memnumber[675 ] = 2'd0;
    assign memnumber[676 ] = 2'd0;
    assign memnumber[677 ] = 2'd0;
    assign memnumber[678 ] = 2'd2;
    assign memnumber[679 ] = 2'd2;
    assign memnumber[680 ] = 2'd1;
    assign memnumber[681 ] = 2'd1;
    assign memnumber[682 ] = 2'd0;
    assign memnumber[683 ] = 2'd0;
    assign memnumber[684 ] = 2'd0;
    assign memnumber[685 ] = 2'd2;
    assign memnumber[686 ] = 2'd2;
    assign memnumber[687 ] = 2'd2;
    assign memnumber[688 ] = 2'd1;
    assign memnumber[689 ] = 2'd1;
    assign memnumber[690 ] = 2'd0;
    assign memnumber[691 ] = 2'd0;
    assign memnumber[692 ] = 2'd0;
    assign memnumber[693 ] = 2'd0;
    assign memnumber[694 ] = 2'd0;
    assign memnumber[695 ] = 2'd0;
    assign memnumber[696 ] = 2'd2;
    assign memnumber[697 ] = 2'd2;
    assign memnumber[698 ] = 2'd2;
    assign memnumber[699 ] = 2'd0;
    assign memnumber[700 ] = 2'd0;
    assign memnumber[701 ] = 2'd0;
    assign memnumber[702 ] = 2'd0;
    assign memnumber[703 ] = 2'd2;
    assign memnumber[704 ] = 2'd2;
    assign memnumber[705 ] = 2'd1;
    assign memnumber[706 ] = 2'd1;
    assign memnumber[707 ] = 2'd1;
    assign memnumber[708 ] = 2'd0;
    assign memnumber[709 ] = 2'd0;
    assign memnumber[710 ] = 2'd0;
    assign memnumber[711 ] = 2'd0;
    assign memnumber[712 ] = 2'd0;
    assign memnumber[713 ] = 2'd1;
    assign memnumber[714 ] = 2'd2;
    assign memnumber[715 ] = 2'd2;
    assign memnumber[716 ] = 2'd0;
    assign memnumber[717 ] = 2'd0;
    assign memnumber[718 ] = 2'd0;
    assign memnumber[719 ] = 2'd0;
    assign memnumber[720 ] = 2'd0;
    assign memnumber[721 ] = 2'd2;
    assign memnumber[722 ] = 2'd2;
    assign memnumber[723 ] = 2'd1;
    assign memnumber[724 ] = 2'd1;
    assign memnumber[725 ] = 2'd0;
    assign memnumber[726 ] = 2'd0;
    assign memnumber[727 ] = 2'd0;
    assign memnumber[728 ] = 2'd0;
    assign memnumber[729 ] = 2'd0;
    assign memnumber[730 ] = 2'd0;
    assign memnumber[731 ] = 2'd0;
    assign memnumber[732 ] = 2'd2;
    assign memnumber[733 ] = 2'd2;
    assign memnumber[734 ] = 2'd2;
    assign memnumber[735 ] = 2'd0;
    assign memnumber[736 ] = 2'd0;
    assign memnumber[737 ] = 2'd0;
    assign memnumber[738 ] = 2'd0;
    assign memnumber[739 ] = 2'd0;
    assign memnumber[740 ] = 2'd0;
    assign memnumber[741 ] = 2'd0;
    assign memnumber[742 ] = 2'd0;
    assign memnumber[743 ] = 2'd0;
    assign memnumber[744 ] = 2'd0;
    assign memnumber[745 ] = 2'd0;
    assign memnumber[746 ] = 2'd2;
    assign memnumber[747 ] = 2'd2;
    assign memnumber[748 ] = 2'd1;
    assign memnumber[749 ] = 2'd0;
    assign memnumber[750 ] = 2'd0;
    assign memnumber[751 ] = 2'd0;
    assign memnumber[752 ] = 2'd0;
    assign memnumber[753 ] = 2'd0;
    assign memnumber[754 ] = 2'd0;
    assign memnumber[755 ] = 2'd0;
    assign memnumber[756 ] = 2'd0;
    assign memnumber[757 ] = 2'd0;
    assign memnumber[758 ] = 2'd2;
    assign memnumber[759 ] = 2'd2;
    assign memnumber[760 ] = 2'd1;
    assign memnumber[761 ] = 2'd1;
    assign memnumber[762 ] = 2'd0;
    assign memnumber[763 ] = 2'd0;
    assign memnumber[764 ] = 2'd0;
    assign memnumber[765 ] = 2'd0;
    assign memnumber[766 ] = 2'd0;
    assign memnumber[767 ] = 2'd0;
    assign memnumber[768 ] = 2'd0;
    assign memnumber[769 ] = 2'd2;
    assign memnumber[770 ] = 2'd2;
    assign memnumber[771 ] = 2'd2;
    assign memnumber[772 ] = 2'd0;
    assign memnumber[773 ] = 2'd0;
    assign memnumber[774 ] = 2'd0;
    assign memnumber[775 ] = 2'd2;
    assign memnumber[776 ] = 2'd2;
    assign memnumber[777 ] = 2'd2;
    assign memnumber[778 ] = 2'd1;
    assign memnumber[779 ] = 2'd0;
    assign memnumber[780 ] = 2'd0;
    assign memnumber[781 ] = 2'd0;
    assign memnumber[782 ] = 2'd0;
    assign memnumber[783 ] = 2'd0;
    assign memnumber[784 ] = 2'd0;
    assign memnumber[785 ] = 2'd0;
    assign memnumber[786 ] = 2'd0;
    assign memnumber[787 ] = 2'd2;
    assign memnumber[788 ] = 2'd2;
    assign memnumber[789 ] = 2'd1;
    assign memnumber[790 ] = 2'd0;
    assign memnumber[791 ] = 2'd0;
    assign memnumber[792 ] = 2'd0;
    assign memnumber[793 ] = 2'd0;
    assign memnumber[794 ] = 2'd0;
    assign memnumber[795 ] = 2'd0;
    assign memnumber[796 ] = 2'd0;
    assign memnumber[797 ] = 2'd0;
    assign memnumber[798 ] = 2'd0;
    assign memnumber[799 ] = 2'd0;
    assign memnumber[800 ] = 2'd0;
    assign memnumber[801 ] = 2'd2;
    assign memnumber[802 ] = 2'd2;
    assign memnumber[803 ] = 2'd2;
    assign memnumber[804 ] = 2'd2;
    assign memnumber[805 ] = 2'd1;
    assign memnumber[806 ] = 2'd0;
    assign memnumber[807 ] = 2'd0;
    assign memnumber[808 ] = 2'd0;
    assign memnumber[809 ] = 2'd0;
    assign memnumber[810 ] = 2'd0;
    assign memnumber[811 ] = 2'd0;
    assign memnumber[812 ] = 2'd0;
    assign memnumber[813 ] = 2'd2;
    assign memnumber[814 ] = 2'd2;
    assign memnumber[815 ] = 2'd1;
    assign memnumber[816 ] = 2'd0;
    assign memnumber[817 ] = 2'd0;
    assign memnumber[818 ] = 2'd0;
    assign memnumber[819 ] = 2'd0;
    assign memnumber[820 ] = 2'd0;
    assign memnumber[821 ] = 2'd0;
    assign memnumber[822 ] = 2'd0;
    assign memnumber[823 ] = 2'd0;
    assign memnumber[824 ] = 2'd0;
    assign memnumber[825 ] = 2'd0;
    assign memnumber[826 ] = 2'd0;
    assign memnumber[827 ] = 2'd0;
    assign memnumber[828 ] = 2'd0;
    assign memnumber[829 ] = 2'd0;
    assign memnumber[830 ] = 2'd0;
    assign memnumber[831 ] = 2'd0;
    assign memnumber[832 ] = 2'd0;
    assign memnumber[833 ] = 2'd0;
    assign memnumber[834 ] = 2'd0;
    assign memnumber[835 ] = 2'd2;
    assign memnumber[836 ] = 2'd2;
    assign memnumber[837 ] = 2'd1;
    assign memnumber[838 ] = 2'd1;
    assign memnumber[839 ] = 2'd0;
    assign memnumber[840 ] = 2'd0;
    assign memnumber[841 ] = 2'd0;
    assign memnumber[842 ] = 2'd0;
    assign memnumber[843 ] = 2'd0;
    assign memnumber[844 ] = 2'd0;
    assign memnumber[845 ] = 2'd0;
    assign memnumber[846 ] = 2'd0;
    assign memnumber[847 ] = 2'd0;
    assign memnumber[848 ] = 2'd0;
    assign memnumber[849 ] = 2'd0;
    assign memnumber[850 ] = 2'd0;
    assign memnumber[851 ] = 2'd0;
    assign memnumber[852 ] = 2'd0;
    assign memnumber[853 ] = 2'd0;
    assign memnumber[854 ] = 2'd0;
    assign memnumber[855 ] = 2'd0;
    assign memnumber[856 ] = 2'd0;
    assign memnumber[857 ] = 2'd0;
    assign memnumber[858 ] = 2'd2;
    assign memnumber[859 ] = 2'd2;
    assign memnumber[860 ] = 2'd1;
    assign memnumber[861 ] = 2'd0;
    assign memnumber[862 ] = 2'd0;
    assign memnumber[863 ] = 2'd0;
    assign memnumber[864 ] = 2'd0;
    assign memnumber[865 ] = 2'd2;
    assign memnumber[866 ] = 2'd2;
    assign memnumber[867 ] = 2'd1;
    assign memnumber[868 ] = 2'd1;
    assign memnumber[869 ] = 2'd0;
    assign memnumber[870 ] = 2'd0;
    assign memnumber[871 ] = 2'd0;
    assign memnumber[872 ] = 2'd0;
    assign memnumber[873 ] = 2'd0;
    assign memnumber[874 ] = 2'd0;
    assign memnumber[875 ] = 2'd0;
    assign memnumber[876 ] = 2'd0;
    assign memnumber[877 ] = 2'd2;
    assign memnumber[878 ] = 2'd2;
    assign memnumber[879 ] = 2'd1;
    assign memnumber[880 ] = 2'd0;
    assign memnumber[881 ] = 2'd0;
    assign memnumber[882 ] = 2'd2;
    assign memnumber[883 ] = 2'd2;
    assign memnumber[884 ] = 2'd2;
    assign memnumber[885 ] = 2'd1;
    assign memnumber[886 ] = 2'd0;
    assign memnumber[887 ] = 2'd0;
    assign memnumber[888 ] = 2'd0;
    assign memnumber[889 ] = 2'd0;
    assign memnumber[890 ] = 2'd0;
    assign memnumber[891 ] = 2'd0;
    assign memnumber[892 ] = 2'd0;
    assign memnumber[893 ] = 2'd0;
    assign memnumber[894 ] = 2'd2;
    assign memnumber[895 ] = 2'd2;
    assign memnumber[896 ] = 2'd2;
    assign memnumber[897 ] = 2'd0;
    assign memnumber[898 ] = 2'd0;
    assign memnumber[899 ] = 2'd0;
    assign memnumber[900 ] = 2'd0;
    assign memnumber[901 ] = 2'd2;
    assign memnumber[902 ] = 2'd2;
    assign memnumber[903 ] = 2'd1;
    assign memnumber[904 ] = 2'd0;
    assign memnumber[905 ] = 2'd0;
    assign memnumber[906 ] = 2'd0;
    assign memnumber[907 ] = 2'd0;
    assign memnumber[908 ] = 2'd0;
    assign memnumber[909 ] = 2'd0;
    assign memnumber[910 ] = 2'd0;
    assign memnumber[911 ] = 2'd0;
    assign memnumber[912 ] = 2'd0;
    assign memnumber[913 ] = 2'd2;
    assign memnumber[914 ] = 2'd2;
    assign memnumber[915 ] = 2'd1;
    assign memnumber[916 ] = 2'd0;
    assign memnumber[917 ] = 2'd0;
    assign memnumber[918 ] = 2'd0;
    assign memnumber[919 ] = 2'd0;
    assign memnumber[920 ] = 2'd0;
    assign memnumber[921 ] = 2'd0;
    assign memnumber[922 ] = 2'd0;
    assign memnumber[923 ] = 2'd0;
    assign memnumber[924 ] = 2'd0;
    assign memnumber[925 ] = 2'd0;
    assign memnumber[926 ] = 2'd2;
    assign memnumber[927 ] = 2'd2;
    assign memnumber[928 ] = 2'd1;
    assign memnumber[929 ] = 2'd0;
    assign memnumber[930 ] = 2'd0;
    assign memnumber[931 ] = 2'd0;
    assign memnumber[932 ] = 2'd0;
    assign memnumber[933 ] = 2'd0;
    assign memnumber[934 ] = 2'd0;
    assign memnumber[935 ] = 2'd0;
    assign memnumber[936 ] = 2'd0;
    assign memnumber[937 ] = 2'd2;
    assign memnumber[938 ] = 2'd2;
    assign memnumber[939 ] = 2'd1;
    assign memnumber[940 ] = 2'd1;
    assign memnumber[941 ] = 2'd0;
    assign memnumber[942 ] = 2'd0;
    assign memnumber[943 ] = 2'd0;
    assign memnumber[944 ] = 2'd0;
    assign memnumber[945 ] = 2'd0;
    assign memnumber[946 ] = 2'd0;
    assign memnumber[947 ] = 2'd0;
    assign memnumber[948 ] = 2'd0;
    assign memnumber[949 ] = 2'd0;
    assign memnumber[950 ] = 2'd2;
    assign memnumber[951 ] = 2'd2;
    assign memnumber[952 ] = 2'd1;
    assign memnumber[953 ] = 2'd0;
    assign memnumber[954 ] = 2'd0;
    assign memnumber[955 ] = 2'd2;
    assign memnumber[956 ] = 2'd2;
    assign memnumber[957 ] = 2'd1;
    assign memnumber[958 ] = 2'd1;
    assign memnumber[959 ] = 2'd0;
    assign memnumber[960 ] = 2'd0;
    assign memnumber[961 ] = 2'd0;
    assign memnumber[962 ] = 2'd0;
    assign memnumber[963 ] = 2'd0;
    assign memnumber[964 ] = 2'd0;
    assign memnumber[965 ] = 2'd0;
    assign memnumber[966 ] = 2'd0;
    assign memnumber[967 ] = 2'd2;
    assign memnumber[968 ] = 2'd2;
    assign memnumber[969 ] = 2'd1;
    assign memnumber[970 ] = 2'd0;
    assign memnumber[971 ] = 2'd0;
    assign memnumber[972 ] = 2'd0;
    assign memnumber[973 ] = 2'd0;
    assign memnumber[974 ] = 2'd0;
    assign memnumber[975 ] = 2'd0;
    assign memnumber[976 ] = 2'd0;
    assign memnumber[977 ] = 2'd0;
    assign memnumber[978 ] = 2'd0;
    assign memnumber[979 ] = 2'd0;
    assign memnumber[980 ] = 2'd0;
    assign memnumber[981 ] = 2'd2;
    assign memnumber[982 ] = 2'd2;
    assign memnumber[983 ] = 2'd2;
    assign memnumber[984 ] = 2'd2;
    assign memnumber[985 ] = 2'd1;
    assign memnumber[986 ] = 2'd0;
    assign memnumber[987 ] = 2'd0;
    assign memnumber[988 ] = 2'd0;
    assign memnumber[989 ] = 2'd0;
    assign memnumber[990 ] = 2'd0;
    assign memnumber[991 ] = 2'd0;
    assign memnumber[992 ] = 2'd0;
    assign memnumber[993 ] = 2'd2;
    assign memnumber[994 ] = 2'd2;
    assign memnumber[995 ] = 2'd1;
    assign memnumber[996 ] = 2'd0;
    assign memnumber[997 ] = 2'd0;
    assign memnumber[998 ] = 2'd0;
    assign memnumber[999 ] = 2'd0;
    assign memnumber[1000] = 2'd0;
    assign memnumber[1001] = 2'd0;
    assign memnumber[1002] = 2'd0;
    assign memnumber[1003] = 2'd0;
    assign memnumber[1004] = 2'd0;
    assign memnumber[1005] = 2'd0;
    assign memnumber[1006] = 2'd0;
    assign memnumber[1007] = 2'd0;
    assign memnumber[1008] = 2'd0;
    assign memnumber[1009] = 2'd0;
    assign memnumber[1010] = 2'd0;
    assign memnumber[1011] = 2'd0;
    assign memnumber[1012] = 2'd0;
    assign memnumber[1013] = 2'd0;
    assign memnumber[1014] = 2'd2;
    assign memnumber[1015] = 2'd2;
    assign memnumber[1016] = 2'd2;
    assign memnumber[1017] = 2'd1;
    assign memnumber[1018] = 2'd0;
    assign memnumber[1019] = 2'd0;
    assign memnumber[1020] = 2'd0;
    assign memnumber[1021] = 2'd0;
    assign memnumber[1022] = 2'd0;
    assign memnumber[1023] = 2'd0;
    assign memnumber[1024] = 2'd0;
    assign memnumber[1025] = 2'd0;
    assign memnumber[1026] = 2'd0;
    assign memnumber[1027] = 2'd0;
    assign memnumber[1028] = 2'd0;
    assign memnumber[1029] = 2'd0;
    assign memnumber[1030] = 2'd0;
    assign memnumber[1031] = 2'd0;
    assign memnumber[1032] = 2'd0;
    assign memnumber[1033] = 2'd0;
    assign memnumber[1034] = 2'd0;
    assign memnumber[1035] = 2'd0;
    assign memnumber[1036] = 2'd0;
    assign memnumber[1037] = 2'd2;
    assign memnumber[1038] = 2'd2;
    assign memnumber[1039] = 2'd1;
    assign memnumber[1040] = 2'd1;
    assign memnumber[1041] = 2'd0;
    assign memnumber[1042] = 2'd0;
    assign memnumber[1043] = 2'd0;
    assign memnumber[1044] = 2'd0;
    assign memnumber[1045] = 2'd2;
    assign memnumber[1046] = 2'd2;
    assign memnumber[1047] = 2'd1;
    assign memnumber[1048] = 2'd0;
    assign memnumber[1049] = 2'd0;
    assign memnumber[1050] = 2'd0;
    assign memnumber[1051] = 2'd0;
    assign memnumber[1052] = 2'd0;
    assign memnumber[1053] = 2'd0;
    assign memnumber[1054] = 2'd0;
    assign memnumber[1055] = 2'd0;
    assign memnumber[1056] = 2'd0;
    assign memnumber[1057] = 2'd2;
    assign memnumber[1058] = 2'd2;
    assign memnumber[1059] = 2'd1;
    assign memnumber[1060] = 2'd0;
    assign memnumber[1061] = 2'd0;
    assign memnumber[1062] = 2'd2;
    assign memnumber[1063] = 2'd2;
    assign memnumber[1064] = 2'd1;
    assign memnumber[1065] = 2'd1;
    assign memnumber[1066] = 2'd0;
    assign memnumber[1067] = 2'd0;
    assign memnumber[1068] = 2'd0;
    assign memnumber[1069] = 2'd0;
    assign memnumber[1070] = 2'd0;
    assign memnumber[1071] = 2'd0;
    assign memnumber[1072] = 2'd0;
    assign memnumber[1073] = 2'd0;
    assign memnumber[1074] = 2'd0;
    assign memnumber[1075] = 2'd2;
    assign memnumber[1076] = 2'd2;
    assign memnumber[1077] = 2'd1;
    assign memnumber[1078] = 2'd0;
    assign memnumber[1079] = 2'd0;
    assign memnumber[1080] = 2'd2;
    assign memnumber[1081] = 2'd2;
    assign memnumber[1082] = 2'd2;
    assign memnumber[1083] = 2'd1;
    assign memnumber[1084] = 2'd0;
    assign memnumber[1085] = 2'd0;
    assign memnumber[1086] = 2'd0;
    assign memnumber[1087] = 2'd0;
    assign memnumber[1088] = 2'd0;
    assign memnumber[1089] = 2'd0;
    assign memnumber[1090] = 2'd0;
    assign memnumber[1091] = 2'd0;
    assign memnumber[1092] = 2'd0;
    assign memnumber[1093] = 2'd2;
    assign memnumber[1094] = 2'd2;
    assign memnumber[1095] = 2'd1;
    assign memnumber[1096] = 2'd0;
    assign memnumber[1097] = 2'd0;
    assign memnumber[1098] = 2'd0;
    assign memnumber[1099] = 2'd0;
    assign memnumber[1100] = 2'd0;
    assign memnumber[1101] = 2'd0;
    assign memnumber[1102] = 2'd0;
    assign memnumber[1103] = 2'd0;
    assign memnumber[1104] = 2'd0;
    assign memnumber[1105] = 2'd0;
    assign memnumber[1106] = 2'd2;
    assign memnumber[1107] = 2'd2;
    assign memnumber[1108] = 2'd1;
    assign memnumber[1109] = 2'd0;
    assign memnumber[1110] = 2'd0;
    assign memnumber[1111] = 2'd0;
    assign memnumber[1112] = 2'd0;
    assign memnumber[1113] = 2'd0;
    assign memnumber[1114] = 2'd0;
    assign memnumber[1115] = 2'd0;
    assign memnumber[1116] = 2'd0;
    assign memnumber[1117] = 2'd2;
    assign memnumber[1118] = 2'd2;
    assign memnumber[1119] = 2'd1;
    assign memnumber[1120] = 2'd0;
    assign memnumber[1121] = 2'd0;
    assign memnumber[1122] = 2'd0;
    assign memnumber[1123] = 2'd0;
    assign memnumber[1124] = 2'd0;
    assign memnumber[1125] = 2'd0;
    assign memnumber[1126] = 2'd0;
    assign memnumber[1127] = 2'd0;
    assign memnumber[1128] = 2'd0;
    assign memnumber[1129] = 2'd0;
    assign memnumber[1130] = 2'd2;
    assign memnumber[1131] = 2'd2;
    assign memnumber[1132] = 2'd1;
    assign memnumber[1133] = 2'd0;
    assign memnumber[1134] = 2'd0;
    assign memnumber[1135] = 2'd0;
    assign memnumber[1136] = 2'd1;
    assign memnumber[1137] = 2'd1;
    assign memnumber[1138] = 2'd0;
    assign memnumber[1139] = 2'd0;
    assign memnumber[1140] = 2'd0;
    assign memnumber[1141] = 2'd0;
    assign memnumber[1142] = 2'd0;
    assign memnumber[1143] = 2'd0;
    assign memnumber[1144] = 2'd0;
    assign memnumber[1145] = 2'd0;
    assign memnumber[1146] = 2'd0;
    assign memnumber[1147] = 2'd2;
    assign memnumber[1148] = 2'd2;
    assign memnumber[1149] = 2'd1;
    assign memnumber[1150] = 2'd0;
    assign memnumber[1151] = 2'd0;
    assign memnumber[1152] = 2'd0;
    assign memnumber[1153] = 2'd0;
    assign memnumber[1154] = 2'd0;
    assign memnumber[1155] = 2'd0;
    assign memnumber[1156] = 2'd0;
    assign memnumber[1157] = 2'd0;
    assign memnumber[1158] = 2'd0;
    assign memnumber[1159] = 2'd0;
    assign memnumber[1160] = 2'd2;
    assign memnumber[1161] = 2'd2;
    assign memnumber[1162] = 2'd1;
    assign memnumber[1163] = 2'd2;
    assign memnumber[1164] = 2'd2;
    assign memnumber[1165] = 2'd1;
    assign memnumber[1166] = 2'd0;
    assign memnumber[1167] = 2'd0;
    assign memnumber[1168] = 2'd0;
    assign memnumber[1169] = 2'd0;
    assign memnumber[1170] = 2'd0;
    assign memnumber[1171] = 2'd0;
    assign memnumber[1172] = 2'd0;
    assign memnumber[1173] = 2'd2;
    assign memnumber[1174] = 2'd2;
    assign memnumber[1175] = 2'd1;
    assign memnumber[1176] = 2'd0;
    assign memnumber[1177] = 2'd0;
    assign memnumber[1178] = 2'd0;
    assign memnumber[1179] = 2'd0;
    assign memnumber[1180] = 2'd0;
    assign memnumber[1181] = 2'd0;
    assign memnumber[1182] = 2'd0;
    assign memnumber[1183] = 2'd0;
    assign memnumber[1184] = 2'd0;
    assign memnumber[1185] = 2'd0;
    assign memnumber[1186] = 2'd0;
    assign memnumber[1187] = 2'd0;
    assign memnumber[1188] = 2'd0;
    assign memnumber[1189] = 2'd0;
    assign memnumber[1190] = 2'd0;
    assign memnumber[1191] = 2'd0;
    assign memnumber[1192] = 2'd0;
    assign memnumber[1193] = 2'd0;
    assign memnumber[1194] = 2'd2;
    assign memnumber[1195] = 2'd2;
    assign memnumber[1196] = 2'd1;
    assign memnumber[1197] = 2'd1;
    assign memnumber[1198] = 2'd0;
    assign memnumber[1199] = 2'd0;
    assign memnumber[1200] = 2'd0;
    assign memnumber[1201] = 2'd0;
    assign memnumber[1202] = 2'd0;
    assign memnumber[1203] = 2'd0;
    assign memnumber[1204] = 2'd0;
    assign memnumber[1205] = 2'd0;
    assign memnumber[1206] = 2'd0;
    assign memnumber[1207] = 2'd0;
    assign memnumber[1208] = 2'd0;
    assign memnumber[1209] = 2'd0;
    assign memnumber[1210] = 2'd0;
    assign memnumber[1211] = 2'd0;
    assign memnumber[1212] = 2'd0;
    assign memnumber[1213] = 2'd0;
    assign memnumber[1214] = 2'd0;
    assign memnumber[1215] = 2'd0;
    assign memnumber[1216] = 2'd2;
    assign memnumber[1217] = 2'd2;
    assign memnumber[1218] = 2'd2;
    assign memnumber[1219] = 2'd1;
    assign memnumber[1220] = 2'd0;
    assign memnumber[1221] = 2'd0;
    assign memnumber[1222] = 2'd0;
    assign memnumber[1223] = 2'd0;
    assign memnumber[1224] = 2'd0;
    assign memnumber[1225] = 2'd2;
    assign memnumber[1226] = 2'd2;
    assign memnumber[1227] = 2'd1;
    assign memnumber[1228] = 2'd0;
    assign memnumber[1229] = 2'd0;
    assign memnumber[1230] = 2'd0;
    assign memnumber[1231] = 2'd0;
    assign memnumber[1232] = 2'd0;
    assign memnumber[1233] = 2'd0;
    assign memnumber[1234] = 2'd0;
    assign memnumber[1235] = 2'd0;
    assign memnumber[1236] = 2'd0;
    assign memnumber[1237] = 2'd2;
    assign memnumber[1238] = 2'd2;
    assign memnumber[1239] = 2'd1;
    assign memnumber[1240] = 2'd0;
    assign memnumber[1241] = 2'd0;
    assign memnumber[1242] = 2'd2;
    assign memnumber[1243] = 2'd2;
    assign memnumber[1244] = 2'd1;
    assign memnumber[1245] = 2'd0;
    assign memnumber[1246] = 2'd0;
    assign memnumber[1247] = 2'd0;
    assign memnumber[1248] = 2'd0;
    assign memnumber[1249] = 2'd0;
    assign memnumber[1250] = 2'd0;
    assign memnumber[1251] = 2'd0;
    assign memnumber[1252] = 2'd0;
    assign memnumber[1253] = 2'd0;
    assign memnumber[1254] = 2'd0;
    assign memnumber[1255] = 2'd2;
    assign memnumber[1256] = 2'd2;
    assign memnumber[1257] = 2'd1;
    assign memnumber[1258] = 2'd0;
    assign memnumber[1259] = 2'd0;
    assign memnumber[1260] = 2'd2;
    assign memnumber[1261] = 2'd2;
    assign memnumber[1262] = 2'd1;
    assign memnumber[1263] = 2'd1;
    assign memnumber[1264] = 2'd0;
    assign memnumber[1265] = 2'd0;
    assign memnumber[1266] = 2'd0;
    assign memnumber[1267] = 2'd0;
    assign memnumber[1268] = 2'd0;
    assign memnumber[1269] = 2'd0;
    assign memnumber[1270] = 2'd0;
    assign memnumber[1271] = 2'd0;
    assign memnumber[1272] = 2'd0;
    assign memnumber[1273] = 2'd0;
    assign memnumber[1274] = 2'd2;
    assign memnumber[1275] = 2'd2;
    assign memnumber[1276] = 2'd0;
    assign memnumber[1277] = 2'd0;
    assign memnumber[1278] = 2'd0;
    assign memnumber[1279] = 2'd0;
    assign memnumber[1280] = 2'd0;
    assign memnumber[1281] = 2'd0;
    assign memnumber[1282] = 2'd0;
    assign memnumber[1283] = 2'd0;
    assign memnumber[1284] = 2'd0;
    assign memnumber[1285] = 2'd0;
    assign memnumber[1286] = 2'd2;
    assign memnumber[1287] = 2'd2;
    assign memnumber[1288] = 2'd1;
    assign memnumber[1289] = 2'd0;
    assign memnumber[1290] = 2'd0;
    assign memnumber[1291] = 2'd0;
    assign memnumber[1292] = 2'd0;
    assign memnumber[1293] = 2'd0;
    assign memnumber[1294] = 2'd0;
    assign memnumber[1295] = 2'd0;
    assign memnumber[1296] = 2'd0;
    assign memnumber[1297] = 2'd0;
    assign memnumber[1298] = 2'd1;
    assign memnumber[1299] = 2'd1;
    assign memnumber[1300] = 2'd0;
    assign memnumber[1301] = 2'd0;
    assign memnumber[1302] = 2'd0;
    assign memnumber[1303] = 2'd0;
    assign memnumber[1304] = 2'd0;
    assign memnumber[1305] = 2'd0;
    assign memnumber[1306] = 2'd0;
    assign memnumber[1307] = 2'd0;
    assign memnumber[1308] = 2'd0;
    assign memnumber[1309] = 2'd0;
    assign memnumber[1310] = 2'd2;
    assign memnumber[1311] = 2'd2;
    assign memnumber[1312] = 2'd1;
    assign memnumber[1313] = 2'd0;
    assign memnumber[1314] = 2'd0;
    assign memnumber[1315] = 2'd0;
    assign memnumber[1316] = 2'd0;
    assign memnumber[1317] = 2'd0;
    assign memnumber[1318] = 2'd0;
    assign memnumber[1319] = 2'd0;
    assign memnumber[1320] = 2'd0;
    assign memnumber[1321] = 2'd0;
    assign memnumber[1322] = 2'd0;
    assign memnumber[1323] = 2'd0;
    assign memnumber[1324] = 2'd0;
    assign memnumber[1325] = 2'd0;
    assign memnumber[1326] = 2'd2;
    assign memnumber[1327] = 2'd2;
    assign memnumber[1328] = 2'd2;
    assign memnumber[1329] = 2'd1;
    assign memnumber[1330] = 2'd0;
    assign memnumber[1331] = 2'd0;
    assign memnumber[1332] = 2'd0;
    assign memnumber[1333] = 2'd0;
    assign memnumber[1334] = 2'd0;
    assign memnumber[1335] = 2'd0;
    assign memnumber[1336] = 2'd0;
    assign memnumber[1337] = 2'd0;
    assign memnumber[1338] = 2'd0;
    assign memnumber[1339] = 2'd2;
    assign memnumber[1340] = 2'd2;
    assign memnumber[1341] = 2'd2;
    assign memnumber[1342] = 2'd1;
    assign memnumber[1343] = 2'd2;
    assign memnumber[1344] = 2'd2;
    assign memnumber[1345] = 2'd1;
    assign memnumber[1346] = 2'd0;
    assign memnumber[1347] = 2'd0;
    assign memnumber[1348] = 2'd0;
    assign memnumber[1349] = 2'd0;
    assign memnumber[1350] = 2'd0;
    assign memnumber[1351] = 2'd0;
    assign memnumber[1352] = 2'd0;
    assign memnumber[1353] = 2'd2;
    assign memnumber[1354] = 2'd2;
    assign memnumber[1355] = 2'd1;
    assign memnumber[1356] = 2'd0;
    assign memnumber[1357] = 2'd0;
    assign memnumber[1358] = 2'd0;
    assign memnumber[1359] = 2'd0;
    assign memnumber[1360] = 2'd0;
    assign memnumber[1361] = 2'd0;
    assign memnumber[1362] = 2'd0;
    assign memnumber[1363] = 2'd0;
    assign memnumber[1364] = 2'd0;
    assign memnumber[1365] = 2'd0;
    assign memnumber[1366] = 2'd0;
    assign memnumber[1367] = 2'd0;
    assign memnumber[1368] = 2'd0;
    assign memnumber[1369] = 2'd0;
    assign memnumber[1370] = 2'd0;
    assign memnumber[1371] = 2'd0;
    assign memnumber[1372] = 2'd0;
    assign memnumber[1373] = 2'd2;
    assign memnumber[1374] = 2'd2;
    assign memnumber[1375] = 2'd1;
    assign memnumber[1376] = 2'd1;
    assign memnumber[1377] = 2'd0;
    assign memnumber[1378] = 2'd0;
    assign memnumber[1379] = 2'd0;
    assign memnumber[1380] = 2'd0;
    assign memnumber[1381] = 2'd0;
    assign memnumber[1382] = 2'd0;
    assign memnumber[1383] = 2'd0;
    assign memnumber[1384] = 2'd0;
    assign memnumber[1385] = 2'd0;
    assign memnumber[1386] = 2'd0;
    assign memnumber[1387] = 2'd0;
    assign memnumber[1388] = 2'd0;
    assign memnumber[1389] = 2'd0;
    assign memnumber[1390] = 2'd0;
    assign memnumber[1391] = 2'd0;
    assign memnumber[1392] = 2'd0;
    assign memnumber[1393] = 2'd0;
    assign memnumber[1394] = 2'd0;
    assign memnumber[1395] = 2'd0;
    assign memnumber[1396] = 2'd2;
    assign memnumber[1397] = 2'd2;
    assign memnumber[1398] = 2'd1;
    assign memnumber[1399] = 2'd1;
    assign memnumber[1400] = 2'd0;
    assign memnumber[1401] = 2'd0;
    assign memnumber[1402] = 2'd0;
    assign memnumber[1403] = 2'd0;
    assign memnumber[1404] = 2'd0;
    assign memnumber[1405] = 2'd0;
    assign memnumber[1406] = 2'd2;
    assign memnumber[1407] = 2'd2;
    assign memnumber[1408] = 2'd0;
    assign memnumber[1409] = 2'd0;
    assign memnumber[1410] = 2'd0;
    assign memnumber[1411] = 2'd0;
    assign memnumber[1412] = 2'd0;
    assign memnumber[1413] = 2'd0;
    assign memnumber[1414] = 2'd0;
    assign memnumber[1415] = 2'd0;
    assign memnumber[1416] = 2'd2;
    assign memnumber[1417] = 2'd2;
    assign memnumber[1418] = 2'd1;
    assign memnumber[1419] = 2'd1;
    assign memnumber[1420] = 2'd0;
    assign memnumber[1421] = 2'd0;
    assign memnumber[1422] = 2'd2;
    assign memnumber[1423] = 2'd2;
    assign memnumber[1424] = 2'd1;
    assign memnumber[1425] = 2'd0;
    assign memnumber[1426] = 2'd0;
    assign memnumber[1427] = 2'd0;
    assign memnumber[1428] = 2'd0;
    assign memnumber[1429] = 2'd0;
    assign memnumber[1430] = 2'd0;
    assign memnumber[1431] = 2'd0;
    assign memnumber[1432] = 2'd0;
    assign memnumber[1433] = 2'd0;
    assign memnumber[1434] = 2'd0;
    assign memnumber[1435] = 2'd2;
    assign memnumber[1436] = 2'd2;
    assign memnumber[1437] = 2'd1;
    assign memnumber[1438] = 2'd0;
    assign memnumber[1439] = 2'd0;
    assign memnumber[1440] = 2'd2;
    assign memnumber[1441] = 2'd2;
    assign memnumber[1442] = 2'd1;
    assign memnumber[1443] = 2'd0;
    assign memnumber[1444] = 2'd0;
    assign memnumber[1445] = 2'd0;
    assign memnumber[1446] = 2'd0;
    assign memnumber[1447] = 2'd0;
    assign memnumber[1448] = 2'd0;
    assign memnumber[1449] = 2'd0;
    assign memnumber[1450] = 2'd0;
    assign memnumber[1451] = 2'd0;
    assign memnumber[1452] = 2'd0;
    assign memnumber[1453] = 2'd0;
    assign memnumber[1454] = 2'd2;
    assign memnumber[1455] = 2'd2;
    assign memnumber[1456] = 2'd1;
    assign memnumber[1457] = 2'd0;
    assign memnumber[1458] = 2'd0;
    assign memnumber[1459] = 2'd0;
    assign memnumber[1460] = 2'd0;
    assign memnumber[1461] = 2'd0;
    assign memnumber[1462] = 2'd0;
    assign memnumber[1463] = 2'd0;
    assign memnumber[1464] = 2'd0;
    assign memnumber[1465] = 2'd0;
    assign memnumber[1466] = 2'd2;
    assign memnumber[1467] = 2'd2;
    assign memnumber[1468] = 2'd1;
    assign memnumber[1469] = 2'd0;
    assign memnumber[1470] = 2'd0;
    assign memnumber[1471] = 2'd0;
    assign memnumber[1472] = 2'd0;
    assign memnumber[1473] = 2'd0;
    assign memnumber[1474] = 2'd0;
    assign memnumber[1475] = 2'd0;
    assign memnumber[1476] = 2'd0;
    assign memnumber[1477] = 2'd0;
    assign memnumber[1478] = 2'd0;
    assign memnumber[1479] = 2'd0;
    assign memnumber[1480] = 2'd0;
    assign memnumber[1481] = 2'd0;
    assign memnumber[1482] = 2'd0;
    assign memnumber[1483] = 2'd0;
    assign memnumber[1484] = 2'd0;
    assign memnumber[1485] = 2'd0;
    assign memnumber[1486] = 2'd0;
    assign memnumber[1487] = 2'd0;
    assign memnumber[1488] = 2'd0;
    assign memnumber[1489] = 2'd0;
    assign memnumber[1490] = 2'd2;
    assign memnumber[1491] = 2'd2;
    assign memnumber[1492] = 2'd1;
    assign memnumber[1493] = 2'd0;
    assign memnumber[1494] = 2'd0;
    assign memnumber[1495] = 2'd0;
    assign memnumber[1496] = 2'd0;
    assign memnumber[1497] = 2'd0;
    assign memnumber[1498] = 2'd0;
    assign memnumber[1499] = 2'd0;
    assign memnumber[1500] = 2'd0;
    assign memnumber[1501] = 2'd0;
    assign memnumber[1502] = 2'd0;
    assign memnumber[1503] = 2'd0;
    assign memnumber[1504] = 2'd2;
    assign memnumber[1505] = 2'd2;
    assign memnumber[1506] = 2'd2;
    assign memnumber[1507] = 2'd2;
    assign memnumber[1508] = 2'd1;
    assign memnumber[1509] = 2'd1;
    assign memnumber[1510] = 2'd0;
    assign memnumber[1511] = 2'd0;
    assign memnumber[1512] = 2'd0;
    assign memnumber[1513] = 2'd0;
    assign memnumber[1514] = 2'd0;
    assign memnumber[1515] = 2'd0;
    assign memnumber[1516] = 2'd0;
    assign memnumber[1517] = 2'd0;
    assign memnumber[1518] = 2'd0;
    assign memnumber[1519] = 2'd2;
    assign memnumber[1520] = 2'd2;
    assign memnumber[1521] = 2'd1;
    assign memnumber[1522] = 2'd1;
    assign memnumber[1523] = 2'd2;
    assign memnumber[1524] = 2'd2;
    assign memnumber[1525] = 2'd1;
    assign memnumber[1526] = 2'd0;
    assign memnumber[1527] = 2'd0;
    assign memnumber[1528] = 2'd0;
    assign memnumber[1529] = 2'd0;
    assign memnumber[1530] = 2'd0;
    assign memnumber[1531] = 2'd0;
    assign memnumber[1532] = 2'd2;
    assign memnumber[1533] = 2'd2;
    assign memnumber[1534] = 2'd2;
    assign memnumber[1535] = 2'd2;
    assign memnumber[1536] = 2'd2;
    assign memnumber[1537] = 2'd2;
    assign memnumber[1538] = 2'd2;
    assign memnumber[1539] = 2'd2;
    assign memnumber[1540] = 2'd0;
    assign memnumber[1541] = 2'd0;
    assign memnumber[1542] = 2'd0;
    assign memnumber[1543] = 2'd0;
    assign memnumber[1544] = 2'd0;
    assign memnumber[1545] = 2'd0;
    assign memnumber[1546] = 2'd0;
    assign memnumber[1547] = 2'd0;
    assign memnumber[1548] = 2'd0;
    assign memnumber[1549] = 2'd0;
    assign memnumber[1550] = 2'd0;
    assign memnumber[1551] = 2'd0;
    assign memnumber[1552] = 2'd2;
    assign memnumber[1553] = 2'd2;
    assign memnumber[1554] = 2'd2;
    assign memnumber[1555] = 2'd1;
    assign memnumber[1556] = 2'd0;
    assign memnumber[1557] = 2'd0;
    assign memnumber[1558] = 2'd0;
    assign memnumber[1559] = 2'd0;
    assign memnumber[1560] = 2'd0;
    assign memnumber[1561] = 2'd0;
    assign memnumber[1562] = 2'd0;
    assign memnumber[1563] = 2'd0;
    assign memnumber[1564] = 2'd0;
    assign memnumber[1565] = 2'd0;
    assign memnumber[1566] = 2'd0;
    assign memnumber[1567] = 2'd0;
    assign memnumber[1568] = 2'd0;
    assign memnumber[1569] = 2'd0;
    assign memnumber[1570] = 2'd0;
    assign memnumber[1571] = 2'd0;
    assign memnumber[1572] = 2'd0;
    assign memnumber[1573] = 2'd0;
    assign memnumber[1574] = 2'd0;
    assign memnumber[1575] = 2'd2;
    assign memnumber[1576] = 2'd2;
    assign memnumber[1577] = 2'd2;
    assign memnumber[1578] = 2'd1;
    assign memnumber[1579] = 2'd0;
    assign memnumber[1580] = 2'd0;
    assign memnumber[1581] = 2'd0;
    assign memnumber[1582] = 2'd0;
    assign memnumber[1583] = 2'd0;
    assign memnumber[1584] = 2'd0;
    assign memnumber[1585] = 2'd0;
    assign memnumber[1586] = 2'd2;
    assign memnumber[1587] = 2'd2;
    assign memnumber[1588] = 2'd2;
    assign memnumber[1589] = 2'd2;
    assign memnumber[1590] = 2'd0;
    assign memnumber[1591] = 2'd0;
    assign memnumber[1592] = 2'd0;
    assign memnumber[1593] = 2'd0;
    assign memnumber[1594] = 2'd0;
    assign memnumber[1595] = 2'd2;
    assign memnumber[1596] = 2'd2;
    assign memnumber[1597] = 2'd2;
    assign memnumber[1598] = 2'd1;
    assign memnumber[1599] = 2'd0;
    assign memnumber[1600] = 2'd0;
    assign memnumber[1601] = 2'd0;
    assign memnumber[1602] = 2'd2;
    assign memnumber[1603] = 2'd2;
    assign memnumber[1604] = 2'd2;
    assign memnumber[1605] = 2'd0;
    assign memnumber[1606] = 2'd0;
    assign memnumber[1607] = 2'd0;
    assign memnumber[1608] = 2'd0;
    assign memnumber[1609] = 2'd0;
    assign memnumber[1610] = 2'd0;
    assign memnumber[1611] = 2'd0;
    assign memnumber[1612] = 2'd0;
    assign memnumber[1613] = 2'd0;
    assign memnumber[1614] = 2'd0;
    assign memnumber[1615] = 2'd2;
    assign memnumber[1616] = 2'd2;
    assign memnumber[1617] = 2'd1;
    assign memnumber[1618] = 2'd0;
    assign memnumber[1619] = 2'd0;
    assign memnumber[1620] = 2'd2;
    assign memnumber[1621] = 2'd2;
    assign memnumber[1622] = 2'd1;
    assign memnumber[1623] = 2'd0;
    assign memnumber[1624] = 2'd0;
    assign memnumber[1625] = 2'd0;
    assign memnumber[1626] = 2'd0;
    assign memnumber[1627] = 2'd0;
    assign memnumber[1628] = 2'd0;
    assign memnumber[1629] = 2'd0;
    assign memnumber[1630] = 2'd0;
    assign memnumber[1631] = 2'd0;
    assign memnumber[1632] = 2'd0;
    assign memnumber[1633] = 2'd0;
    assign memnumber[1634] = 2'd2;
    assign memnumber[1635] = 2'd2;
    assign memnumber[1636] = 2'd1;
    assign memnumber[1637] = 2'd0;
    assign memnumber[1638] = 2'd0;
    assign memnumber[1639] = 2'd0;
    assign memnumber[1640] = 2'd0;
    assign memnumber[1641] = 2'd0;
    assign memnumber[1642] = 2'd0;
    assign memnumber[1643] = 2'd0;
    assign memnumber[1644] = 2'd0;
    assign memnumber[1645] = 2'd0;
    assign memnumber[1646] = 2'd2;
    assign memnumber[1647] = 2'd2;
    assign memnumber[1648] = 2'd1;
    assign memnumber[1649] = 2'd0;
    assign memnumber[1650] = 2'd0;
    assign memnumber[1651] = 2'd0;
    assign memnumber[1652] = 2'd0;
    assign memnumber[1653] = 2'd0;
    assign memnumber[1654] = 2'd0;
    assign memnumber[1655] = 2'd0;
    assign memnumber[1656] = 2'd0;
    assign memnumber[1657] = 2'd0;
    assign memnumber[1658] = 2'd0;
    assign memnumber[1659] = 2'd0;
    assign memnumber[1660] = 2'd0;
    assign memnumber[1661] = 2'd0;
    assign memnumber[1662] = 2'd0;
    assign memnumber[1663] = 2'd0;
    assign memnumber[1664] = 2'd0;
    assign memnumber[1665] = 2'd0;
    assign memnumber[1666] = 2'd0;
    assign memnumber[1667] = 2'd0;
    assign memnumber[1668] = 2'd0;
    assign memnumber[1669] = 2'd2;
    assign memnumber[1670] = 2'd2;
    assign memnumber[1671] = 2'd1;
    assign memnumber[1672] = 2'd1;
    assign memnumber[1673] = 2'd0;
    assign memnumber[1674] = 2'd0;
    assign memnumber[1675] = 2'd0;
    assign memnumber[1676] = 2'd0;
    assign memnumber[1677] = 2'd0;
    assign memnumber[1678] = 2'd0;
    assign memnumber[1679] = 2'd0;
    assign memnumber[1680] = 2'd0;
    assign memnumber[1681] = 2'd2;
    assign memnumber[1682] = 2'd2;
    assign memnumber[1683] = 2'd2;
    assign memnumber[1684] = 2'd2;
    assign memnumber[1685] = 2'd2;
    assign memnumber[1686] = 2'd2;
    assign memnumber[1687] = 2'd1;
    assign memnumber[1688] = 2'd1;
    assign memnumber[1689] = 2'd0;
    assign memnumber[1690] = 2'd0;
    assign memnumber[1691] = 2'd0;
    assign memnumber[1692] = 2'd0;
    assign memnumber[1693] = 2'd0;
    assign memnumber[1694] = 2'd0;
    assign memnumber[1695] = 2'd0;
    assign memnumber[1696] = 2'd0;
    assign memnumber[1697] = 2'd0;
    assign memnumber[1698] = 2'd2;
    assign memnumber[1699] = 2'd2;
    assign memnumber[1700] = 2'd1;
    assign memnumber[1701] = 2'd1;
    assign memnumber[1702] = 2'd0;
    assign memnumber[1703] = 2'd2;
    assign memnumber[1704] = 2'd2;
    assign memnumber[1705] = 2'd1;
    assign memnumber[1706] = 2'd0;
    assign memnumber[1707] = 2'd0;
    assign memnumber[1708] = 2'd0;
    assign memnumber[1709] = 2'd0;
    assign memnumber[1710] = 2'd0;
    assign memnumber[1711] = 2'd0;
    assign memnumber[1712] = 2'd2;
    assign memnumber[1713] = 2'd2;
    assign memnumber[1714] = 2'd2;
    assign memnumber[1715] = 2'd2;
    assign memnumber[1716] = 2'd2;
    assign memnumber[1717] = 2'd2;
    assign memnumber[1718] = 2'd2;
    assign memnumber[1719] = 2'd2;
    assign memnumber[1720] = 2'd2;
    assign memnumber[1721] = 2'd2;
    assign memnumber[1722] = 2'd0;
    assign memnumber[1723] = 2'd0;
    assign memnumber[1724] = 2'd0;
    assign memnumber[1725] = 2'd0;
    assign memnumber[1726] = 2'd0;
    assign memnumber[1727] = 2'd0;
    assign memnumber[1728] = 2'd0;
    assign memnumber[1729] = 2'd0;
    assign memnumber[1730] = 2'd0;
    assign memnumber[1731] = 2'd0;
    assign memnumber[1732] = 2'd2;
    assign memnumber[1733] = 2'd2;
    assign memnumber[1734] = 2'd1;
    assign memnumber[1735] = 2'd1;
    assign memnumber[1736] = 2'd0;
    assign memnumber[1737] = 2'd0;
    assign memnumber[1738] = 2'd0;
    assign memnumber[1739] = 2'd0;
    assign memnumber[1740] = 2'd0;
    assign memnumber[1741] = 2'd0;
    assign memnumber[1742] = 2'd0;
    assign memnumber[1743] = 2'd0;
    assign memnumber[1744] = 2'd0;
    assign memnumber[1745] = 2'd0;
    assign memnumber[1746] = 2'd0;
    assign memnumber[1747] = 2'd0;
    assign memnumber[1748] = 2'd0;
    assign memnumber[1749] = 2'd0;
    assign memnumber[1750] = 2'd0;
    assign memnumber[1751] = 2'd0;
    assign memnumber[1752] = 2'd0;
    assign memnumber[1753] = 2'd0;
    assign memnumber[1754] = 2'd0;
    assign memnumber[1755] = 2'd2;
    assign memnumber[1756] = 2'd2;
    assign memnumber[1757] = 2'd1;
    assign memnumber[1758] = 2'd1;
    assign memnumber[1759] = 2'd0;
    assign memnumber[1760] = 2'd0;
    assign memnumber[1761] = 2'd0;
    assign memnumber[1762] = 2'd0;
    assign memnumber[1763] = 2'd0;
    assign memnumber[1764] = 2'd0;
    assign memnumber[1765] = 2'd0;
    assign memnumber[1766] = 2'd0;
    assign memnumber[1767] = 2'd1;
    assign memnumber[1768] = 2'd2;
    assign memnumber[1769] = 2'd2;
    assign memnumber[1770] = 2'd2;
    assign memnumber[1771] = 2'd2;
    assign memnumber[1772] = 2'd2;
    assign memnumber[1773] = 2'd2;
    assign memnumber[1774] = 2'd2;
    assign memnumber[1775] = 2'd2;
    assign memnumber[1776] = 2'd1;
    assign memnumber[1777] = 2'd1;
    assign memnumber[1778] = 2'd1;
    assign memnumber[1779] = 2'd0;
    assign memnumber[1780] = 2'd0;
    assign memnumber[1781] = 2'd0;
    assign memnumber[1782] = 2'd0;
    assign memnumber[1783] = 2'd2;
    assign memnumber[1784] = 2'd2;
    assign memnumber[1785] = 2'd2;
    assign memnumber[1786] = 2'd0;
    assign memnumber[1787] = 2'd0;
    assign memnumber[1788] = 2'd0;
    assign memnumber[1789] = 2'd0;
    assign memnumber[1790] = 2'd0;
    assign memnumber[1791] = 2'd0;
    assign memnumber[1792] = 2'd0;
    assign memnumber[1793] = 2'd0;
    assign memnumber[1794] = 2'd2;
    assign memnumber[1795] = 2'd2;
    assign memnumber[1796] = 2'd1;
    assign memnumber[1797] = 2'd1;
    assign memnumber[1798] = 2'd0;
    assign memnumber[1799] = 2'd0;
    assign memnumber[1800] = 2'd2;
    assign memnumber[1801] = 2'd2;
    assign memnumber[1802] = 2'd1;
    assign memnumber[1803] = 2'd0;
    assign memnumber[1804] = 2'd0;
    assign memnumber[1805] = 2'd0;
    assign memnumber[1806] = 2'd0;
    assign memnumber[1807] = 2'd0;
    assign memnumber[1808] = 2'd0;
    assign memnumber[1809] = 2'd0;
    assign memnumber[1810] = 2'd0;
    assign memnumber[1811] = 2'd0;
    assign memnumber[1812] = 2'd0;
    assign memnumber[1813] = 2'd0;
    assign memnumber[1814] = 2'd2;
    assign memnumber[1815] = 2'd2;
    assign memnumber[1816] = 2'd1;
    assign memnumber[1817] = 2'd0;
    assign memnumber[1818] = 2'd0;
    assign memnumber[1819] = 2'd0;
    assign memnumber[1820] = 2'd0;
    assign memnumber[1821] = 2'd0;
    assign memnumber[1822] = 2'd0;
    assign memnumber[1823] = 2'd0;
    assign memnumber[1824] = 2'd0;
    assign memnumber[1825] = 2'd0;
    assign memnumber[1826] = 2'd2;
    assign memnumber[1827] = 2'd2;
    assign memnumber[1828] = 2'd1;
    assign memnumber[1829] = 2'd0;
    assign memnumber[1830] = 2'd0;
    assign memnumber[1831] = 2'd0;
    assign memnumber[1832] = 2'd0;
    assign memnumber[1833] = 2'd0;
    assign memnumber[1834] = 2'd0;
    assign memnumber[1835] = 2'd0;
    assign memnumber[1836] = 2'd0;
    assign memnumber[1837] = 2'd0;
    assign memnumber[1838] = 2'd0;
    assign memnumber[1839] = 2'd0;
    assign memnumber[1840] = 2'd0;
    assign memnumber[1841] = 2'd0;
    assign memnumber[1842] = 2'd0;
    assign memnumber[1843] = 2'd0;
    assign memnumber[1844] = 2'd0;
    assign memnumber[1845] = 2'd0;
    assign memnumber[1846] = 2'd0;
    assign memnumber[1847] = 2'd0;
    assign memnumber[1848] = 2'd2;
    assign memnumber[1849] = 2'd2;
    assign memnumber[1850] = 2'd2;
    assign memnumber[1851] = 2'd1;
    assign memnumber[1852] = 2'd0;
    assign memnumber[1853] = 2'd0;
    assign memnumber[1854] = 2'd0;
    assign memnumber[1855] = 2'd0;
    assign memnumber[1856] = 2'd0;
    assign memnumber[1857] = 2'd0;
    assign memnumber[1858] = 2'd0;
    assign memnumber[1859] = 2'd0;
    assign memnumber[1860] = 2'd0;
    assign memnumber[1861] = 2'd2;
    assign memnumber[1862] = 2'd2;
    assign memnumber[1863] = 2'd2;
    assign memnumber[1864] = 2'd2;
    assign memnumber[1865] = 2'd2;
    assign memnumber[1866] = 2'd2;
    assign memnumber[1867] = 2'd1;
    assign memnumber[1868] = 2'd0;
    assign memnumber[1869] = 2'd0;
    assign memnumber[1870] = 2'd0;
    assign memnumber[1871] = 2'd0;
    assign memnumber[1872] = 2'd0;
    assign memnumber[1873] = 2'd0;
    assign memnumber[1874] = 2'd0;
    assign memnumber[1875] = 2'd0;
    assign memnumber[1876] = 2'd0;
    assign memnumber[1877] = 2'd2;
    assign memnumber[1878] = 2'd2;
    assign memnumber[1879] = 2'd1;
    assign memnumber[1880] = 2'd1;
    assign memnumber[1881] = 2'd0;
    assign memnumber[1882] = 2'd0;
    assign memnumber[1883] = 2'd2;
    assign memnumber[1884] = 2'd2;
    assign memnumber[1885] = 2'd1;
    assign memnumber[1886] = 2'd0;
    assign memnumber[1887] = 2'd0;
    assign memnumber[1888] = 2'd0;
    assign memnumber[1889] = 2'd0;
    assign memnumber[1890] = 2'd0;
    assign memnumber[1891] = 2'd0;
    assign memnumber[1892] = 2'd2;
    assign memnumber[1893] = 2'd2;
    assign memnumber[1894] = 2'd1;
    assign memnumber[1895] = 2'd1;
    assign memnumber[1896] = 2'd1;
    assign memnumber[1897] = 2'd1;
    assign memnumber[1898] = 2'd1;
    assign memnumber[1899] = 2'd1;
    assign memnumber[1900] = 2'd2;
    assign memnumber[1901] = 2'd2;
    assign memnumber[1902] = 2'd2;
    assign memnumber[1903] = 2'd0;
    assign memnumber[1904] = 2'd0;
    assign memnumber[1905] = 2'd0;
    assign memnumber[1906] = 2'd0;
    assign memnumber[1907] = 2'd0;
    assign memnumber[1908] = 2'd0;
    assign memnumber[1909] = 2'd0;
    assign memnumber[1910] = 2'd0;
    assign memnumber[1911] = 2'd2;
    assign memnumber[1912] = 2'd2;
    assign memnumber[1913] = 2'd2;
    assign memnumber[1914] = 2'd2;
    assign memnumber[1915] = 2'd2;
    assign memnumber[1916] = 2'd2;
    assign memnumber[1917] = 2'd2;
    assign memnumber[1918] = 2'd2;
    assign memnumber[1919] = 2'd0;
    assign memnumber[1920] = 2'd0;
    assign memnumber[1921] = 2'd0;
    assign memnumber[1922] = 2'd0;
    assign memnumber[1923] = 2'd0;
    assign memnumber[1924] = 2'd0;
    assign memnumber[1925] = 2'd0;
    assign memnumber[1926] = 2'd0;
    assign memnumber[1927] = 2'd0;
    assign memnumber[1928] = 2'd0;
    assign memnumber[1929] = 2'd0;
    assign memnumber[1930] = 2'd0;
    assign memnumber[1931] = 2'd0;
    assign memnumber[1932] = 2'd0;
    assign memnumber[1933] = 2'd0;
    assign memnumber[1934] = 2'd2;
    assign memnumber[1935] = 2'd2;
    assign memnumber[1936] = 2'd2;
    assign memnumber[1937] = 2'd1;
    assign memnumber[1938] = 2'd0;
    assign memnumber[1939] = 2'd0;
    assign memnumber[1940] = 2'd0;
    assign memnumber[1941] = 2'd0;
    assign memnumber[1942] = 2'd0;
    assign memnumber[1943] = 2'd0;
    assign memnumber[1944] = 2'd0;
    assign memnumber[1945] = 2'd0;
    assign memnumber[1946] = 2'd0;
    assign memnumber[1947] = 2'd2;
    assign memnumber[1948] = 2'd2;
    assign memnumber[1949] = 2'd2;
    assign memnumber[1950] = 2'd2;
    assign memnumber[1951] = 2'd2;
    assign memnumber[1952] = 2'd2;
    assign memnumber[1953] = 2'd2;
    assign memnumber[1954] = 2'd2;
    assign memnumber[1955] = 2'd2;
    assign memnumber[1956] = 2'd2;
    assign memnumber[1957] = 2'd0;
    assign memnumber[1958] = 2'd0;
    assign memnumber[1959] = 2'd0;
    assign memnumber[1960] = 2'd0;
    assign memnumber[1961] = 2'd0;
    assign memnumber[1962] = 2'd0;
    assign memnumber[1963] = 2'd0;
    assign memnumber[1964] = 2'd2;
    assign memnumber[1965] = 2'd2;
    assign memnumber[1966] = 2'd2;
    assign memnumber[1967] = 2'd0;
    assign memnumber[1968] = 2'd0;
    assign memnumber[1969] = 2'd0;
    assign memnumber[1970] = 2'd0;
    assign memnumber[1971] = 2'd0;
    assign memnumber[1972] = 2'd0;
    assign memnumber[1973] = 2'd2;
    assign memnumber[1974] = 2'd2;
    assign memnumber[1975] = 2'd2;
    assign memnumber[1976] = 2'd1;
    assign memnumber[1977] = 2'd0;
    assign memnumber[1978] = 2'd0;
    assign memnumber[1979] = 2'd0;
    assign memnumber[1980] = 2'd2;
    assign memnumber[1981] = 2'd2;
    assign memnumber[1982] = 2'd1;
    assign memnumber[1983] = 2'd0;
    assign memnumber[1984] = 2'd0;
    assign memnumber[1985] = 2'd0;
    assign memnumber[1986] = 2'd0;
    assign memnumber[1987] = 2'd0;
    assign memnumber[1988] = 2'd0;
    assign memnumber[1989] = 2'd0;
    assign memnumber[1990] = 2'd0;
    assign memnumber[1991] = 2'd0;
    assign memnumber[1992] = 2'd0;
    assign memnumber[1993] = 2'd0;
    assign memnumber[1994] = 2'd2;
    assign memnumber[1995] = 2'd2;
    assign memnumber[1996] = 2'd1;
    assign memnumber[1997] = 2'd0;
    assign memnumber[1998] = 2'd0;
    assign memnumber[1999] = 2'd0;
    assign memnumber[2000] = 2'd0;
    assign memnumber[2001] = 2'd0;
    assign memnumber[2002] = 2'd0;
    assign memnumber[2003] = 2'd0;
    assign memnumber[2004] = 2'd0;
    assign memnumber[2005] = 2'd0;
    assign memnumber[2006] = 2'd2;
    assign memnumber[2007] = 2'd2;
    assign memnumber[2008] = 2'd1;
    assign memnumber[2009] = 2'd0;
    assign memnumber[2010] = 2'd0;
    assign memnumber[2011] = 2'd0;
    assign memnumber[2012] = 2'd0;
    assign memnumber[2013] = 2'd0;
    assign memnumber[2014] = 2'd0;
    assign memnumber[2015] = 2'd0;
    assign memnumber[2016] = 2'd0;
    assign memnumber[2017] = 2'd0;
    assign memnumber[2018] = 2'd0;
    assign memnumber[2019] = 2'd0;
    assign memnumber[2020] = 2'd0;
    assign memnumber[2021] = 2'd0;
    assign memnumber[2022] = 2'd0;
    assign memnumber[2023] = 2'd0;
    assign memnumber[2024] = 2'd0;
    assign memnumber[2025] = 2'd0;
    assign memnumber[2026] = 2'd0;
    assign memnumber[2027] = 2'd0;
    assign memnumber[2028] = 2'd2;
    assign memnumber[2029] = 2'd2;
    assign memnumber[2030] = 2'd1;
    assign memnumber[2031] = 2'd1;
    assign memnumber[2032] = 2'd0;
    assign memnumber[2033] = 2'd0;
    assign memnumber[2034] = 2'd0;
    assign memnumber[2035] = 2'd0;
    assign memnumber[2036] = 2'd0;
    assign memnumber[2037] = 2'd0;
    assign memnumber[2038] = 2'd0;
    assign memnumber[2039] = 2'd0;
    assign memnumber[2040] = 2'd0;
    assign memnumber[2041] = 2'd0;
    assign memnumber[2042] = 2'd1;
    assign memnumber[2043] = 2'd1;
    assign memnumber[2044] = 2'd2;
    assign memnumber[2045] = 2'd2;
    assign memnumber[2046] = 2'd2;
    assign memnumber[2047] = 2'd2;
    assign memnumber[2048] = 2'd2;
    assign memnumber[2049] = 2'd0;
    assign memnumber[2050] = 2'd0;
    assign memnumber[2051] = 2'd0;
    assign memnumber[2052] = 2'd0;
    assign memnumber[2053] = 2'd0;
    assign memnumber[2054] = 2'd0;
    assign memnumber[2055] = 2'd0;
    assign memnumber[2056] = 2'd0;
    assign memnumber[2057] = 2'd2;
    assign memnumber[2058] = 2'd2;
    assign memnumber[2059] = 2'd1;
    assign memnumber[2060] = 2'd0;
    assign memnumber[2061] = 2'd0;
    assign memnumber[2062] = 2'd0;
    assign memnumber[2063] = 2'd2;
    assign memnumber[2064] = 2'd2;
    assign memnumber[2065] = 2'd1;
    assign memnumber[2066] = 2'd0;
    assign memnumber[2067] = 2'd0;
    assign memnumber[2068] = 2'd0;
    assign memnumber[2069] = 2'd0;
    assign memnumber[2070] = 2'd0;
    assign memnumber[2071] = 2'd0;
    assign memnumber[2072] = 2'd0;
    assign memnumber[2073] = 2'd1;
    assign memnumber[2074] = 2'd1;
    assign memnumber[2075] = 2'd0;
    assign memnumber[2076] = 2'd0;
    assign memnumber[2077] = 2'd0;
    assign memnumber[2078] = 2'd0;
    assign memnumber[2079] = 2'd0;
    assign memnumber[2080] = 2'd0;
    assign memnumber[2081] = 2'd1;
    assign memnumber[2082] = 2'd2;
    assign memnumber[2083] = 2'd2;
    assign memnumber[2084] = 2'd0;
    assign memnumber[2085] = 2'd0;
    assign memnumber[2086] = 2'd0;
    assign memnumber[2087] = 2'd0;
    assign memnumber[2088] = 2'd0;
    assign memnumber[2089] = 2'd0;
    assign memnumber[2090] = 2'd2;
    assign memnumber[2091] = 2'd2;
    assign memnumber[2092] = 2'd2;
    assign memnumber[2093] = 2'd2;
    assign memnumber[2094] = 2'd2;
    assign memnumber[2095] = 2'd2;
    assign memnumber[2096] = 2'd2;
    assign memnumber[2097] = 2'd2;
    assign memnumber[2098] = 2'd2;
    assign memnumber[2099] = 2'd2;
    assign memnumber[2100] = 2'd0;
    assign memnumber[2101] = 2'd0;
    assign memnumber[2102] = 2'd0;
    assign memnumber[2103] = 2'd0;
    assign memnumber[2104] = 2'd0;
    assign memnumber[2105] = 2'd0;
    assign memnumber[2106] = 2'd0;
    assign memnumber[2107] = 2'd0;
    assign memnumber[2108] = 2'd0;
    assign memnumber[2109] = 2'd0;
    assign memnumber[2110] = 2'd0;
    assign memnumber[2111] = 2'd0;
    assign memnumber[2112] = 2'd0;
    assign memnumber[2113] = 2'd0;
    assign memnumber[2114] = 2'd2;
    assign memnumber[2115] = 2'd2;
    assign memnumber[2116] = 2'd1;
    assign memnumber[2117] = 2'd1;
    assign memnumber[2118] = 2'd0;
    assign memnumber[2119] = 2'd0;
    assign memnumber[2120] = 2'd0;
    assign memnumber[2121] = 2'd0;
    assign memnumber[2122] = 2'd0;
    assign memnumber[2123] = 2'd0;
    assign memnumber[2124] = 2'd0;
    assign memnumber[2125] = 2'd0;
    assign memnumber[2126] = 2'd2;
    assign memnumber[2127] = 2'd2;
    assign memnumber[2128] = 2'd2;
    assign memnumber[2129] = 2'd1;
    assign memnumber[2130] = 2'd1;
    assign memnumber[2131] = 2'd1;
    assign memnumber[2132] = 2'd1;
    assign memnumber[2133] = 2'd1;
    assign memnumber[2134] = 2'd1;
    assign memnumber[2135] = 2'd2;
    assign memnumber[2136] = 2'd2;
    assign memnumber[2137] = 2'd2;
    assign memnumber[2138] = 2'd0;
    assign memnumber[2139] = 2'd0;
    assign memnumber[2140] = 2'd0;
    assign memnumber[2141] = 2'd0;
    assign memnumber[2142] = 2'd0;
    assign memnumber[2143] = 2'd0;
    assign memnumber[2144] = 2'd0;
    assign memnumber[2145] = 2'd2;
    assign memnumber[2146] = 2'd2;
    assign memnumber[2147] = 2'd2;
    assign memnumber[2148] = 2'd2;
    assign memnumber[2149] = 2'd2;
    assign memnumber[2150] = 2'd2;
    assign memnumber[2151] = 2'd2;
    assign memnumber[2152] = 2'd2;
    assign memnumber[2153] = 2'd2;
    assign memnumber[2154] = 2'd2;
    assign memnumber[2155] = 2'd1;
    assign memnumber[2156] = 2'd1;
    assign memnumber[2157] = 2'd0;
    assign memnumber[2158] = 2'd0;
    assign memnumber[2159] = 2'd0;
    assign memnumber[2160] = 2'd2;
    assign memnumber[2161] = 2'd2;
    assign memnumber[2162] = 2'd1;
    assign memnumber[2163] = 2'd0;
    assign memnumber[2164] = 2'd0;
    assign memnumber[2165] = 2'd0;
    assign memnumber[2166] = 2'd0;
    assign memnumber[2167] = 2'd0;
    assign memnumber[2168] = 2'd0;
    assign memnumber[2169] = 2'd0;
    assign memnumber[2170] = 2'd0;
    assign memnumber[2171] = 2'd0;
    assign memnumber[2172] = 2'd0;
    assign memnumber[2173] = 2'd0;
    assign memnumber[2174] = 2'd2;
    assign memnumber[2175] = 2'd2;
    assign memnumber[2176] = 2'd1;
    assign memnumber[2177] = 2'd0;
    assign memnumber[2178] = 2'd0;
    assign memnumber[2179] = 2'd0;
    assign memnumber[2180] = 2'd0;
    assign memnumber[2181] = 2'd0;
    assign memnumber[2182] = 2'd0;
    assign memnumber[2183] = 2'd0;
    assign memnumber[2184] = 2'd0;
    assign memnumber[2185] = 2'd0;
    assign memnumber[2186] = 2'd2;
    assign memnumber[2187] = 2'd2;
    assign memnumber[2188] = 2'd1;
    assign memnumber[2189] = 2'd0;
    assign memnumber[2190] = 2'd0;
    assign memnumber[2191] = 2'd0;
    assign memnumber[2192] = 2'd0;
    assign memnumber[2193] = 2'd0;
    assign memnumber[2194] = 2'd0;
    assign memnumber[2195] = 2'd0;
    assign memnumber[2196] = 2'd0;
    assign memnumber[2197] = 2'd0;
    assign memnumber[2198] = 2'd0;
    assign memnumber[2199] = 2'd0;
    assign memnumber[2200] = 2'd0;
    assign memnumber[2201] = 2'd0;
    assign memnumber[2202] = 2'd0;
    assign memnumber[2203] = 2'd0;
    assign memnumber[2204] = 2'd0;
    assign memnumber[2205] = 2'd0;
    assign memnumber[2206] = 2'd0;
    assign memnumber[2207] = 2'd2;
    assign memnumber[2208] = 2'd2;
    assign memnumber[2209] = 2'd1;
    assign memnumber[2210] = 2'd1;
    assign memnumber[2211] = 2'd0;
    assign memnumber[2212] = 2'd0;
    assign memnumber[2213] = 2'd0;
    assign memnumber[2214] = 2'd0;
    assign memnumber[2215] = 2'd0;
    assign memnumber[2216] = 2'd0;
    assign memnumber[2217] = 2'd0;
    assign memnumber[2218] = 2'd0;
    assign memnumber[2219] = 2'd0;
    assign memnumber[2220] = 2'd0;
    assign memnumber[2221] = 2'd0;
    assign memnumber[2222] = 2'd0;
    assign memnumber[2223] = 2'd0;
    assign memnumber[2224] = 2'd0;
    assign memnumber[2225] = 2'd1;
    assign memnumber[2226] = 2'd2;
    assign memnumber[2227] = 2'd2;
    assign memnumber[2228] = 2'd2;
    assign memnumber[2229] = 2'd1;
    assign memnumber[2230] = 2'd0;
    assign memnumber[2231] = 2'd0;
    assign memnumber[2232] = 2'd0;
    assign memnumber[2233] = 2'd0;
    assign memnumber[2234] = 2'd0;
    assign memnumber[2235] = 2'd0;
    assign memnumber[2236] = 2'd2;
    assign memnumber[2237] = 2'd2;
    assign memnumber[2238] = 2'd1;
    assign memnumber[2239] = 2'd1;
    assign memnumber[2240] = 2'd0;
    assign memnumber[2241] = 2'd0;
    assign memnumber[2242] = 2'd0;
    assign memnumber[2243] = 2'd2;
    assign memnumber[2244] = 2'd2;
    assign memnumber[2245] = 2'd1;
    assign memnumber[2246] = 2'd0;
    assign memnumber[2247] = 2'd0;
    assign memnumber[2248] = 2'd0;
    assign memnumber[2249] = 2'd0;
    assign memnumber[2250] = 2'd0;
    assign memnumber[2251] = 2'd0;
    assign memnumber[2252] = 2'd0;
    assign memnumber[2253] = 2'd0;
    assign memnumber[2254] = 2'd0;
    assign memnumber[2255] = 2'd0;
    assign memnumber[2256] = 2'd0;
    assign memnumber[2257] = 2'd0;
    assign memnumber[2258] = 2'd0;
    assign memnumber[2259] = 2'd0;
    assign memnumber[2260] = 2'd0;
    assign memnumber[2261] = 2'd0;
    assign memnumber[2262] = 2'd2;
    assign memnumber[2263] = 2'd2;
    assign memnumber[2264] = 2'd2;
    assign memnumber[2265] = 2'd0;
    assign memnumber[2266] = 2'd0;
    assign memnumber[2267] = 2'd0;
    assign memnumber[2268] = 2'd0;
    assign memnumber[2269] = 2'd0;
    assign memnumber[2270] = 2'd2;
    assign memnumber[2271] = 2'd2;
    assign memnumber[2272] = 2'd2;
    assign memnumber[2273] = 2'd1;
    assign memnumber[2274] = 2'd1;
    assign memnumber[2275] = 2'd1;
    assign memnumber[2276] = 2'd1;
    assign memnumber[2277] = 2'd1;
    assign memnumber[2278] = 2'd2;
    assign memnumber[2279] = 2'd2;
    assign memnumber[2280] = 2'd2;
    assign memnumber[2281] = 2'd2;
    assign memnumber[2282] = 2'd0;
    assign memnumber[2283] = 2'd0;
    assign memnumber[2284] = 2'd0;
    assign memnumber[2285] = 2'd0;
    assign memnumber[2286] = 2'd0;
    assign memnumber[2287] = 2'd0;
    assign memnumber[2288] = 2'd0;
    assign memnumber[2289] = 2'd0;
    assign memnumber[2290] = 2'd0;
    assign memnumber[2291] = 2'd0;
    assign memnumber[2292] = 2'd0;
    assign memnumber[2293] = 2'd2;
    assign memnumber[2294] = 2'd2;
    assign memnumber[2295] = 2'd1;
    assign memnumber[2296] = 2'd1;
    assign memnumber[2297] = 2'd0;
    assign memnumber[2298] = 2'd0;
    assign memnumber[2299] = 2'd0;
    assign memnumber[2300] = 2'd0;
    assign memnumber[2301] = 2'd0;
    assign memnumber[2302] = 2'd0;
    assign memnumber[2303] = 2'd0;
    assign memnumber[2304] = 2'd0;
    assign memnumber[2305] = 2'd2;
    assign memnumber[2306] = 2'd2;
    assign memnumber[2307] = 2'd2;
    assign memnumber[2308] = 2'd1;
    assign memnumber[2309] = 2'd1;
    assign memnumber[2310] = 2'd0;
    assign memnumber[2311] = 2'd0;
    assign memnumber[2312] = 2'd0;
    assign memnumber[2313] = 2'd0;
    assign memnumber[2314] = 2'd0;
    assign memnumber[2315] = 2'd0;
    assign memnumber[2316] = 2'd2;
    assign memnumber[2317] = 2'd2;
    assign memnumber[2318] = 2'd2;
    assign memnumber[2319] = 2'd0;
    assign memnumber[2320] = 2'd0;
    assign memnumber[2321] = 2'd0;
    assign memnumber[2322] = 2'd0;
    assign memnumber[2323] = 2'd0;
    assign memnumber[2324] = 2'd0;
    assign memnumber[2325] = 2'd0;
    assign memnumber[2326] = 2'd1;
    assign memnumber[2327] = 2'd2;
    assign memnumber[2328] = 2'd2;
    assign memnumber[2329] = 2'd2;
    assign memnumber[2330] = 2'd2;
    assign memnumber[2331] = 2'd2;
    assign memnumber[2332] = 2'd2;
    assign memnumber[2333] = 2'd2;
    assign memnumber[2334] = 2'd2;
    assign memnumber[2335] = 2'd1;
    assign memnumber[2336] = 2'd0;
    assign memnumber[2337] = 2'd0;
    assign memnumber[2338] = 2'd0;
    assign memnumber[2339] = 2'd0;
    assign memnumber[2340] = 2'd2;
    assign memnumber[2341] = 2'd2;
    assign memnumber[2342] = 2'd1;
    assign memnumber[2343] = 2'd0;
    assign memnumber[2344] = 2'd0;
    assign memnumber[2345] = 2'd0;
    assign memnumber[2346] = 2'd0;
    assign memnumber[2347] = 2'd0;
    assign memnumber[2348] = 2'd0;
    assign memnumber[2349] = 2'd0;
    assign memnumber[2350] = 2'd0;
    assign memnumber[2351] = 2'd0;
    assign memnumber[2352] = 2'd0;
    assign memnumber[2353] = 2'd0;
    assign memnumber[2354] = 2'd2;
    assign memnumber[2355] = 2'd2;
    assign memnumber[2356] = 2'd1;
    assign memnumber[2357] = 2'd0;
    assign memnumber[2358] = 2'd0;
    assign memnumber[2359] = 2'd0;
    assign memnumber[2360] = 2'd0;
    assign memnumber[2361] = 2'd0;
    assign memnumber[2362] = 2'd0;
    assign memnumber[2363] = 2'd0;
    assign memnumber[2364] = 2'd0;
    assign memnumber[2365] = 2'd0;
    assign memnumber[2366] = 2'd2;
    assign memnumber[2367] = 2'd2;
    assign memnumber[2368] = 2'd1;
    assign memnumber[2369] = 2'd0;
    assign memnumber[2370] = 2'd0;
    assign memnumber[2371] = 2'd0;
    assign memnumber[2372] = 2'd0;
    assign memnumber[2373] = 2'd0;
    assign memnumber[2374] = 2'd0;
    assign memnumber[2375] = 2'd0;
    assign memnumber[2376] = 2'd0;
    assign memnumber[2377] = 2'd0;
    assign memnumber[2378] = 2'd0;
    assign memnumber[2379] = 2'd0;
    assign memnumber[2380] = 2'd0;
    assign memnumber[2381] = 2'd0;
    assign memnumber[2382] = 2'd0;
    assign memnumber[2383] = 2'd0;
    assign memnumber[2384] = 2'd0;
    assign memnumber[2385] = 2'd0;
    assign memnumber[2386] = 2'd2;
    assign memnumber[2387] = 2'd2;
    assign memnumber[2388] = 2'd1;
    assign memnumber[2389] = 2'd1;
    assign memnumber[2390] = 2'd0;
    assign memnumber[2391] = 2'd0;
    assign memnumber[2392] = 2'd0;
    assign memnumber[2393] = 2'd0;
    assign memnumber[2394] = 2'd0;
    assign memnumber[2395] = 2'd0;
    assign memnumber[2396] = 2'd0;
    assign memnumber[2397] = 2'd0;
    assign memnumber[2398] = 2'd0;
    assign memnumber[2399] = 2'd0;
    assign memnumber[2400] = 2'd0;
    assign memnumber[2401] = 2'd0;
    assign memnumber[2402] = 2'd0;
    assign memnumber[2403] = 2'd0;
    assign memnumber[2404] = 2'd0;
    assign memnumber[2405] = 2'd0;
    assign memnumber[2406] = 2'd0;
    assign memnumber[2407] = 2'd2;
    assign memnumber[2408] = 2'd2;
    assign memnumber[2409] = 2'd2;
    assign memnumber[2410] = 2'd0;
    assign memnumber[2411] = 2'd0;
    assign memnumber[2412] = 2'd0;
    assign memnumber[2413] = 2'd0;
    assign memnumber[2414] = 2'd0;
    assign memnumber[2415] = 2'd2;
    assign memnumber[2416] = 2'd2;
    assign memnumber[2417] = 2'd1;
    assign memnumber[2418] = 2'd1;
    assign memnumber[2419] = 2'd0;
    assign memnumber[2420] = 2'd0;
    assign memnumber[2421] = 2'd0;
    assign memnumber[2422] = 2'd0;
    assign memnumber[2423] = 2'd2;
    assign memnumber[2424] = 2'd2;
    assign memnumber[2425] = 2'd1;
    assign memnumber[2426] = 2'd0;
    assign memnumber[2427] = 2'd0;
    assign memnumber[2428] = 2'd0;
    assign memnumber[2429] = 2'd0;
    assign memnumber[2430] = 2'd0;
    assign memnumber[2431] = 2'd0;
    assign memnumber[2432] = 2'd0;
    assign memnumber[2433] = 2'd0;
    assign memnumber[2434] = 2'd0;
    assign memnumber[2435] = 2'd0;
    assign memnumber[2436] = 2'd0;
    assign memnumber[2437] = 2'd0;
    assign memnumber[2438] = 2'd0;
    assign memnumber[2439] = 2'd0;
    assign memnumber[2440] = 2'd0;
    assign memnumber[2441] = 2'd0;
    assign memnumber[2442] = 2'd0;
    assign memnumber[2443] = 2'd2;
    assign memnumber[2444] = 2'd2;
    assign memnumber[2445] = 2'd1;
    assign memnumber[2446] = 2'd0;
    assign memnumber[2447] = 2'd0;
    assign memnumber[2448] = 2'd0;
    assign memnumber[2449] = 2'd0;
    assign memnumber[2450] = 2'd2;
    assign memnumber[2451] = 2'd2;
    assign memnumber[2452] = 2'd1;
    assign memnumber[2453] = 2'd1;
    assign memnumber[2454] = 2'd0;
    assign memnumber[2455] = 2'd0;
    assign memnumber[2456] = 2'd0;
    assign memnumber[2457] = 2'd0;
    assign memnumber[2458] = 2'd0;
    assign memnumber[2459] = 2'd1;
    assign memnumber[2460] = 2'd2;
    assign memnumber[2461] = 2'd2;
    assign memnumber[2462] = 2'd1;
    assign memnumber[2463] = 2'd0;
    assign memnumber[2464] = 2'd0;
    assign memnumber[2465] = 2'd0;
    assign memnumber[2466] = 2'd0;
    assign memnumber[2467] = 2'd0;
    assign memnumber[2468] = 2'd0;
    assign memnumber[2469] = 2'd0;
    assign memnumber[2470] = 2'd0;
    assign memnumber[2471] = 2'd0;
    assign memnumber[2472] = 2'd0;
    assign memnumber[2473] = 2'd2;
    assign memnumber[2474] = 2'd2;
    assign memnumber[2475] = 2'd1;
    assign memnumber[2476] = 2'd0;
    assign memnumber[2477] = 2'd0;
    assign memnumber[2478] = 2'd0;
    assign memnumber[2479] = 2'd0;
    assign memnumber[2480] = 2'd0;
    assign memnumber[2481] = 2'd0;
    assign memnumber[2482] = 2'd0;
    assign memnumber[2483] = 2'd0;
    assign memnumber[2484] = 2'd0;
    assign memnumber[2485] = 2'd2;
    assign memnumber[2486] = 2'd2;
    assign memnumber[2487] = 2'd1;
    assign memnumber[2488] = 2'd1;
    assign memnumber[2489] = 2'd0;
    assign memnumber[2490] = 2'd0;
    assign memnumber[2491] = 2'd0;
    assign memnumber[2492] = 2'd0;
    assign memnumber[2493] = 2'd0;
    assign memnumber[2494] = 2'd0;
    assign memnumber[2495] = 2'd0;
    assign memnumber[2496] = 2'd0;
    assign memnumber[2497] = 2'd2;
    assign memnumber[2498] = 2'd2;
    assign memnumber[2499] = 2'd2;
    assign memnumber[2500] = 2'd0;
    assign memnumber[2501] = 2'd0;
    assign memnumber[2502] = 2'd0;
    assign memnumber[2503] = 2'd0;
    assign memnumber[2504] = 2'd0;
    assign memnumber[2505] = 2'd0;
    assign memnumber[2506] = 2'd0;
    assign memnumber[2507] = 2'd0;
    assign memnumber[2508] = 2'd1;
    assign memnumber[2509] = 2'd1;
    assign memnumber[2510] = 2'd1;
    assign memnumber[2511] = 2'd1;
    assign memnumber[2512] = 2'd2;
    assign memnumber[2513] = 2'd2;
    assign memnumber[2514] = 2'd1;
    assign memnumber[2515] = 2'd1;
    assign memnumber[2516] = 2'd0;
    assign memnumber[2517] = 2'd0;
    assign memnumber[2518] = 2'd0;
    assign memnumber[2519] = 2'd0;
    assign memnumber[2520] = 2'd2;
    assign memnumber[2521] = 2'd2;
    assign memnumber[2522] = 2'd1;
    assign memnumber[2523] = 2'd0;
    assign memnumber[2524] = 2'd0;
    assign memnumber[2525] = 2'd0;
    assign memnumber[2526] = 2'd0;
    assign memnumber[2527] = 2'd0;
    assign memnumber[2528] = 2'd0;
    assign memnumber[2529] = 2'd0;
    assign memnumber[2530] = 2'd0;
    assign memnumber[2531] = 2'd0;
    assign memnumber[2532] = 2'd0;
    assign memnumber[2533] = 2'd0;
    assign memnumber[2534] = 2'd2;
    assign memnumber[2535] = 2'd2;
    assign memnumber[2536] = 2'd1;
    assign memnumber[2537] = 2'd0;
    assign memnumber[2538] = 2'd0;
    assign memnumber[2539] = 2'd0;
    assign memnumber[2540] = 2'd0;
    assign memnumber[2541] = 2'd0;
    assign memnumber[2542] = 2'd0;
    assign memnumber[2543] = 2'd0;
    assign memnumber[2544] = 2'd0;
    assign memnumber[2545] = 2'd0;
    assign memnumber[2546] = 2'd2;
    assign memnumber[2547] = 2'd2;
    assign memnumber[2548] = 2'd1;
    assign memnumber[2549] = 2'd0;
    assign memnumber[2550] = 2'd0;
    assign memnumber[2551] = 2'd0;
    assign memnumber[2552] = 2'd0;
    assign memnumber[2553] = 2'd0;
    assign memnumber[2554] = 2'd0;
    assign memnumber[2555] = 2'd0;
    assign memnumber[2556] = 2'd0;
    assign memnumber[2557] = 2'd0;
    assign memnumber[2558] = 2'd0;
    assign memnumber[2559] = 2'd0;
    assign memnumber[2560] = 2'd0;
    assign memnumber[2561] = 2'd0;
    assign memnumber[2562] = 2'd0;
    assign memnumber[2563] = 2'd0;
    assign memnumber[2564] = 2'd0;
    assign memnumber[2565] = 2'd2;
    assign memnumber[2566] = 2'd2;
    assign memnumber[2567] = 2'd1;
    assign memnumber[2568] = 2'd1;
    assign memnumber[2569] = 2'd0;
    assign memnumber[2570] = 2'd0;
    assign memnumber[2571] = 2'd0;
    assign memnumber[2572] = 2'd0;
    assign memnumber[2573] = 2'd0;
    assign memnumber[2574] = 2'd0;
    assign memnumber[2575] = 2'd0;
    assign memnumber[2576] = 2'd0;
    assign memnumber[2577] = 2'd0;
    assign memnumber[2578] = 2'd0;
    assign memnumber[2579] = 2'd0;
    assign memnumber[2580] = 2'd0;
    assign memnumber[2581] = 2'd0;
    assign memnumber[2582] = 2'd0;
    assign memnumber[2583] = 2'd0;
    assign memnumber[2584] = 2'd0;
    assign memnumber[2585] = 2'd0;
    assign memnumber[2586] = 2'd0;
    assign memnumber[2587] = 2'd0;
    assign memnumber[2588] = 2'd2;
    assign memnumber[2589] = 2'd2;
    assign memnumber[2590] = 2'd1;
    assign memnumber[2591] = 2'd0;
    assign memnumber[2592] = 2'd0;
    assign memnumber[2593] = 2'd0;
    assign memnumber[2594] = 2'd2;
    assign memnumber[2595] = 2'd2;
    assign memnumber[2596] = 2'd2;
    assign memnumber[2597] = 2'd1;
    assign memnumber[2598] = 2'd0;
    assign memnumber[2599] = 2'd0;
    assign memnumber[2600] = 2'd0;
    assign memnumber[2601] = 2'd0;
    assign memnumber[2602] = 2'd0;
    assign memnumber[2603] = 2'd2;
    assign memnumber[2604] = 2'd2;
    assign memnumber[2605] = 2'd1;
    assign memnumber[2606] = 2'd0;
    assign memnumber[2607] = 2'd0;
    assign memnumber[2608] = 2'd0;
    assign memnumber[2609] = 2'd0;
    assign memnumber[2610] = 2'd0;
    assign memnumber[2611] = 2'd0;
    assign memnumber[2612] = 2'd0;
    assign memnumber[2613] = 2'd0;
    assign memnumber[2614] = 2'd0;
    assign memnumber[2615] = 2'd0;
    assign memnumber[2616] = 2'd0;
    assign memnumber[2617] = 2'd0;
    assign memnumber[2618] = 2'd0;
    assign memnumber[2619] = 2'd0;
    assign memnumber[2620] = 2'd0;
    assign memnumber[2621] = 2'd0;
    assign memnumber[2622] = 2'd0;
    assign memnumber[2623] = 2'd2;
    assign memnumber[2624] = 2'd2;
    assign memnumber[2625] = 2'd1;
    assign memnumber[2626] = 2'd0;
    assign memnumber[2627] = 2'd0;
    assign memnumber[2628] = 2'd0;
    assign memnumber[2629] = 2'd2;
    assign memnumber[2630] = 2'd2;
    assign memnumber[2631] = 2'd1;
    assign memnumber[2632] = 2'd1;
    assign memnumber[2633] = 2'd0;
    assign memnumber[2634] = 2'd0;
    assign memnumber[2635] = 2'd0;
    assign memnumber[2636] = 2'd0;
    assign memnumber[2637] = 2'd0;
    assign memnumber[2638] = 2'd0;
    assign memnumber[2639] = 2'd0;
    assign memnumber[2640] = 2'd2;
    assign memnumber[2641] = 2'd2;
    assign memnumber[2642] = 2'd2;
    assign memnumber[2643] = 2'd0;
    assign memnumber[2644] = 2'd0;
    assign memnumber[2645] = 2'd0;
    assign memnumber[2646] = 2'd0;
    assign memnumber[2647] = 2'd0;
    assign memnumber[2648] = 2'd0;
    assign memnumber[2649] = 2'd0;
    assign memnumber[2650] = 2'd0;
    assign memnumber[2651] = 2'd0;
    assign memnumber[2652] = 2'd2;
    assign memnumber[2653] = 2'd2;
    assign memnumber[2654] = 2'd1;
    assign memnumber[2655] = 2'd1;
    assign memnumber[2656] = 2'd0;
    assign memnumber[2657] = 2'd0;
    assign memnumber[2658] = 2'd0;
    assign memnumber[2659] = 2'd0;
    assign memnumber[2660] = 2'd0;
    assign memnumber[2661] = 2'd0;
    assign memnumber[2662] = 2'd0;
    assign memnumber[2663] = 2'd0;
    assign memnumber[2664] = 2'd2;
    assign memnumber[2665] = 2'd2;
    assign memnumber[2666] = 2'd1;
    assign memnumber[2667] = 2'd1;
    assign memnumber[2668] = 2'd0;
    assign memnumber[2669] = 2'd0;
    assign memnumber[2670] = 2'd0;
    assign memnumber[2671] = 2'd0;
    assign memnumber[2672] = 2'd0;
    assign memnumber[2673] = 2'd0;
    assign memnumber[2674] = 2'd0;
    assign memnumber[2675] = 2'd0;
    assign memnumber[2676] = 2'd0;
    assign memnumber[2677] = 2'd0;
    assign memnumber[2678] = 2'd2;
    assign memnumber[2679] = 2'd2;
    assign memnumber[2680] = 2'd1;
    assign memnumber[2681] = 2'd0;
    assign memnumber[2682] = 2'd0;
    assign memnumber[2683] = 2'd0;
    assign memnumber[2684] = 2'd0;
    assign memnumber[2685] = 2'd0;
    assign memnumber[2686] = 2'd0;
    assign memnumber[2687] = 2'd0;
    assign memnumber[2688] = 2'd0;
    assign memnumber[2689] = 2'd0;
    assign memnumber[2690] = 2'd0;
    assign memnumber[2691] = 2'd2;
    assign memnumber[2692] = 2'd2;
    assign memnumber[2693] = 2'd1;
    assign memnumber[2694] = 2'd1;
    assign memnumber[2695] = 2'd0;
    assign memnumber[2696] = 2'd0;
    assign memnumber[2697] = 2'd0;
    assign memnumber[2698] = 2'd0;
    assign memnumber[2699] = 2'd0;
    assign memnumber[2700] = 2'd2;
    assign memnumber[2701] = 2'd2;
    assign memnumber[2702] = 2'd1;
    assign memnumber[2703] = 2'd0;
    assign memnumber[2704] = 2'd0;
    assign memnumber[2705] = 2'd0;
    assign memnumber[2706] = 2'd0;
    assign memnumber[2707] = 2'd0;
    assign memnumber[2708] = 2'd0;
    assign memnumber[2709] = 2'd0;
    assign memnumber[2710] = 2'd0;
    assign memnumber[2711] = 2'd0;
    assign memnumber[2712] = 2'd0;
    assign memnumber[2713] = 2'd0;
    assign memnumber[2714] = 2'd2;
    assign memnumber[2715] = 2'd2;
    assign memnumber[2716] = 2'd1;
    assign memnumber[2717] = 2'd0;
    assign memnumber[2718] = 2'd0;
    assign memnumber[2719] = 2'd0;
    assign memnumber[2720] = 2'd0;
    assign memnumber[2721] = 2'd0;
    assign memnumber[2722] = 2'd0;
    assign memnumber[2723] = 2'd0;
    assign memnumber[2724] = 2'd0;
    assign memnumber[2725] = 2'd0;
    assign memnumber[2726] = 2'd2;
    assign memnumber[2727] = 2'd2;
    assign memnumber[2728] = 2'd1;
    assign memnumber[2729] = 2'd0;
    assign memnumber[2730] = 2'd0;
    assign memnumber[2731] = 2'd0;
    assign memnumber[2732] = 2'd0;
    assign memnumber[2733] = 2'd0;
    assign memnumber[2734] = 2'd0;
    assign memnumber[2735] = 2'd0;
    assign memnumber[2736] = 2'd0;
    assign memnumber[2737] = 2'd0;
    assign memnumber[2738] = 2'd0;
    assign memnumber[2739] = 2'd0;
    assign memnumber[2740] = 2'd0;
    assign memnumber[2741] = 2'd0;
    assign memnumber[2742] = 2'd0;
    assign memnumber[2743] = 2'd0;
    assign memnumber[2744] = 2'd2;
    assign memnumber[2745] = 2'd2;
    assign memnumber[2746] = 2'd1;
    assign memnumber[2747] = 2'd1;
    assign memnumber[2748] = 2'd0;
    assign memnumber[2749] = 2'd0;
    assign memnumber[2750] = 2'd0;
    assign memnumber[2751] = 2'd0;
    assign memnumber[2752] = 2'd0;
    assign memnumber[2753] = 2'd0;
    assign memnumber[2754] = 2'd0;
    assign memnumber[2755] = 2'd0;
    assign memnumber[2756] = 2'd0;
    assign memnumber[2757] = 2'd0;
    assign memnumber[2758] = 2'd0;
    assign memnumber[2759] = 2'd0;
    assign memnumber[2760] = 2'd0;
    assign memnumber[2761] = 2'd0;
    assign memnumber[2762] = 2'd0;
    assign memnumber[2763] = 2'd0;
    assign memnumber[2764] = 2'd0;
    assign memnumber[2765] = 2'd0;
    assign memnumber[2766] = 2'd0;
    assign memnumber[2767] = 2'd0;
    assign memnumber[2768] = 2'd2;
    assign memnumber[2769] = 2'd2;
    assign memnumber[2770] = 2'd1;
    assign memnumber[2771] = 2'd0;
    assign memnumber[2772] = 2'd0;
    assign memnumber[2773] = 2'd0;
    assign memnumber[2774] = 2'd2;
    assign memnumber[2775] = 2'd2;
    assign memnumber[2776] = 2'd1;
    assign memnumber[2777] = 2'd1;
    assign memnumber[2778] = 2'd0;
    assign memnumber[2779] = 2'd0;
    assign memnumber[2780] = 2'd0;
    assign memnumber[2781] = 2'd0;
    assign memnumber[2782] = 2'd0;
    assign memnumber[2783] = 2'd2;
    assign memnumber[2784] = 2'd2;
    assign memnumber[2785] = 2'd1;
    assign memnumber[2786] = 2'd0;
    assign memnumber[2787] = 2'd0;
    assign memnumber[2788] = 2'd0;
    assign memnumber[2789] = 2'd0;
    assign memnumber[2790] = 2'd0;
    assign memnumber[2791] = 2'd0;
    assign memnumber[2792] = 2'd0;
    assign memnumber[2793] = 2'd0;
    assign memnumber[2794] = 2'd0;
    assign memnumber[2795] = 2'd0;
    assign memnumber[2796] = 2'd0;
    assign memnumber[2797] = 2'd0;
    assign memnumber[2798] = 2'd0;
    assign memnumber[2799] = 2'd0;
    assign memnumber[2800] = 2'd0;
    assign memnumber[2801] = 2'd0;
    assign memnumber[2802] = 2'd0;
    assign memnumber[2803] = 2'd2;
    assign memnumber[2804] = 2'd2;
    assign memnumber[2805] = 2'd1;
    assign memnumber[2806] = 2'd0;
    assign memnumber[2807] = 2'd0;
    assign memnumber[2808] = 2'd0;
    assign memnumber[2809] = 2'd2;
    assign memnumber[2810] = 2'd2;
    assign memnumber[2811] = 2'd1;
    assign memnumber[2812] = 2'd0;
    assign memnumber[2813] = 2'd0;
    assign memnumber[2814] = 2'd0;
    assign memnumber[2815] = 2'd0;
    assign memnumber[2816] = 2'd0;
    assign memnumber[2817] = 2'd0;
    assign memnumber[2818] = 2'd0;
    assign memnumber[2819] = 2'd0;
    assign memnumber[2820] = 2'd0;
    assign memnumber[2821] = 2'd2;
    assign memnumber[2822] = 2'd2;
    assign memnumber[2823] = 2'd1;
    assign memnumber[2824] = 2'd0;
    assign memnumber[2825] = 2'd0;
    assign memnumber[2826] = 2'd0;
    assign memnumber[2827] = 2'd0;
    assign memnumber[2828] = 2'd0;
    assign memnumber[2829] = 2'd0;
    assign memnumber[2830] = 2'd0;
    assign memnumber[2831] = 2'd0;
    assign memnumber[2832] = 2'd2;
    assign memnumber[2833] = 2'd2;
    assign memnumber[2834] = 2'd1;
    assign memnumber[2835] = 2'd0;
    assign memnumber[2836] = 2'd0;
    assign memnumber[2837] = 2'd0;
    assign memnumber[2838] = 2'd0;
    assign memnumber[2839] = 2'd0;
    assign memnumber[2840] = 2'd0;
    assign memnumber[2841] = 2'd0;
    assign memnumber[2842] = 2'd0;
    assign memnumber[2843] = 2'd0;
    assign memnumber[2844] = 2'd2;
    assign memnumber[2845] = 2'd2;
    assign memnumber[2846] = 2'd1;
    assign memnumber[2847] = 2'd0;
    assign memnumber[2848] = 2'd0;
    assign memnumber[2849] = 2'd0;
    assign memnumber[2850] = 2'd0;
    assign memnumber[2851] = 2'd0;
    assign memnumber[2852] = 2'd0;
    assign memnumber[2853] = 2'd0;
    assign memnumber[2854] = 2'd0;
    assign memnumber[2855] = 2'd0;
    assign memnumber[2856] = 2'd0;
    assign memnumber[2857] = 2'd0;
    assign memnumber[2858] = 2'd2;
    assign memnumber[2859] = 2'd2;
    assign memnumber[2860] = 2'd1;
    assign memnumber[2861] = 2'd0;
    assign memnumber[2862] = 2'd0;
    assign memnumber[2863] = 2'd0;
    assign memnumber[2864] = 2'd0;
    assign memnumber[2865] = 2'd0;
    assign memnumber[2866] = 2'd0;
    assign memnumber[2867] = 2'd0;
    assign memnumber[2868] = 2'd0;
    assign memnumber[2869] = 2'd0;
    assign memnumber[2870] = 2'd2;
    assign memnumber[2871] = 2'd2;
    assign memnumber[2872] = 2'd2;
    assign memnumber[2873] = 2'd1;
    assign memnumber[2874] = 2'd0;
    assign memnumber[2875] = 2'd0;
    assign memnumber[2876] = 2'd0;
    assign memnumber[2877] = 2'd0;
    assign memnumber[2878] = 2'd0;
    assign memnumber[2879] = 2'd0;
    assign memnumber[2880] = 2'd2;
    assign memnumber[2881] = 2'd2;
    assign memnumber[2882] = 2'd2;
    assign memnumber[2883] = 2'd0;
    assign memnumber[2884] = 2'd0;
    assign memnumber[2885] = 2'd0;
    assign memnumber[2886] = 2'd0;
    assign memnumber[2887] = 2'd0;
    assign memnumber[2888] = 2'd0;
    assign memnumber[2889] = 2'd0;
    assign memnumber[2890] = 2'd0;
    assign memnumber[2891] = 2'd0;
    assign memnumber[2892] = 2'd0;
    assign memnumber[2893] = 2'd2;
    assign memnumber[2894] = 2'd2;
    assign memnumber[2895] = 2'd1;
    assign memnumber[2896] = 2'd1;
    assign memnumber[2897] = 2'd0;
    assign memnumber[2898] = 2'd0;
    assign memnumber[2899] = 2'd0;
    assign memnumber[2900] = 2'd0;
    assign memnumber[2901] = 2'd0;
    assign memnumber[2902] = 2'd0;
    assign memnumber[2903] = 2'd0;
    assign memnumber[2904] = 2'd0;
    assign memnumber[2905] = 2'd0;
    assign memnumber[2906] = 2'd2;
    assign memnumber[2907] = 2'd2;
    assign memnumber[2908] = 2'd1;
    assign memnumber[2909] = 2'd0;
    assign memnumber[2910] = 2'd0;
    assign memnumber[2911] = 2'd0;
    assign memnumber[2912] = 2'd0;
    assign memnumber[2913] = 2'd0;
    assign memnumber[2914] = 2'd0;
    assign memnumber[2915] = 2'd0;
    assign memnumber[2916] = 2'd0;
    assign memnumber[2917] = 2'd0;
    assign memnumber[2918] = 2'd0;
    assign memnumber[2919] = 2'd0;
    assign memnumber[2920] = 2'd0;
    assign memnumber[2921] = 2'd0;
    assign memnumber[2922] = 2'd0;
    assign memnumber[2923] = 2'd2;
    assign memnumber[2924] = 2'd2;
    assign memnumber[2925] = 2'd1;
    assign memnumber[2926] = 2'd1;
    assign memnumber[2927] = 2'd0;
    assign memnumber[2928] = 2'd0;
    assign memnumber[2929] = 2'd0;
    assign memnumber[2930] = 2'd0;
    assign memnumber[2931] = 2'd0;
    assign memnumber[2932] = 2'd0;
    assign memnumber[2933] = 2'd0;
    assign memnumber[2934] = 2'd2;
    assign memnumber[2935] = 2'd2;
    assign memnumber[2936] = 2'd0;
    assign memnumber[2937] = 2'd0;
    assign memnumber[2938] = 2'd0;
    assign memnumber[2939] = 2'd0;
    assign memnumber[2940] = 2'd0;
    assign memnumber[2941] = 2'd0;
    assign memnumber[2942] = 2'd0;
    assign memnumber[2943] = 2'd0;
    assign memnumber[2944] = 2'd0;
    assign memnumber[2945] = 2'd0;
    assign memnumber[2946] = 2'd0;
    assign memnumber[2947] = 2'd0;
    assign memnumber[2948] = 2'd2;
    assign memnumber[2949] = 2'd2;
    assign memnumber[2950] = 2'd1;
    assign memnumber[2951] = 2'd0;
    assign memnumber[2952] = 2'd0;
    assign memnumber[2953] = 2'd2;
    assign memnumber[2954] = 2'd2;
    assign memnumber[2955] = 2'd2;
    assign memnumber[2956] = 2'd2;
    assign memnumber[2957] = 2'd2;
    assign memnumber[2958] = 2'd2;
    assign memnumber[2959] = 2'd2;
    assign memnumber[2960] = 2'd2;
    assign memnumber[2961] = 2'd2;
    assign memnumber[2962] = 2'd2;
    assign memnumber[2963] = 2'd2;
    assign memnumber[2964] = 2'd2;
    assign memnumber[2965] = 2'd2;
    assign memnumber[2966] = 2'd2;
    assign memnumber[2967] = 2'd2;
    assign memnumber[2968] = 2'd0;
    assign memnumber[2969] = 2'd0;
    assign memnumber[2970] = 2'd0;
    assign memnumber[2971] = 2'd0;
    assign memnumber[2972] = 2'd0;
    assign memnumber[2973] = 2'd0;
    assign memnumber[2974] = 2'd0;
    assign memnumber[2975] = 2'd0;
    assign memnumber[2976] = 2'd0;
    assign memnumber[2977] = 2'd0;
    assign memnumber[2978] = 2'd0;
    assign memnumber[2979] = 2'd0;
    assign memnumber[2980] = 2'd0;
    assign memnumber[2981] = 2'd0;
    assign memnumber[2982] = 2'd0;
    assign memnumber[2983] = 2'd2;
    assign memnumber[2984] = 2'd2;
    assign memnumber[2985] = 2'd1;
    assign memnumber[2986] = 2'd0;
    assign memnumber[2987] = 2'd0;
    assign memnumber[2988] = 2'd0;
    assign memnumber[2989] = 2'd2;
    assign memnumber[2990] = 2'd2;
    assign memnumber[2991] = 2'd1;
    assign memnumber[2992] = 2'd0;
    assign memnumber[2993] = 2'd0;
    assign memnumber[2994] = 2'd0;
    assign memnumber[2995] = 2'd0;
    assign memnumber[2996] = 2'd0;
    assign memnumber[2997] = 2'd0;
    assign memnumber[2998] = 2'd0;
    assign memnumber[2999] = 2'd0;
    assign memnumber[3000] = 2'd0;
    assign memnumber[3001] = 2'd2;
    assign memnumber[3002] = 2'd2;
    assign memnumber[3003] = 2'd1;
    assign memnumber[3004] = 2'd0;
    assign memnumber[3005] = 2'd0;
    assign memnumber[3006] = 2'd0;
    assign memnumber[3007] = 2'd0;
    assign memnumber[3008] = 2'd0;
    assign memnumber[3009] = 2'd0;
    assign memnumber[3010] = 2'd0;
    assign memnumber[3011] = 2'd2;
    assign memnumber[3012] = 2'd2;
    assign memnumber[3013] = 2'd1;
    assign memnumber[3014] = 2'd1;
    assign memnumber[3015] = 2'd0;
    assign memnumber[3016] = 2'd0;
    assign memnumber[3017] = 2'd0;
    assign memnumber[3018] = 2'd0;
    assign memnumber[3019] = 2'd0;
    assign memnumber[3020] = 2'd0;
    assign memnumber[3021] = 2'd0;
    assign memnumber[3022] = 2'd0;
    assign memnumber[3023] = 2'd0;
    assign memnumber[3024] = 2'd2;
    assign memnumber[3025] = 2'd2;
    assign memnumber[3026] = 2'd1;
    assign memnumber[3027] = 2'd0;
    assign memnumber[3028] = 2'd0;
    assign memnumber[3029] = 2'd0;
    assign memnumber[3030] = 2'd0;
    assign memnumber[3031] = 2'd0;
    assign memnumber[3032] = 2'd0;
    assign memnumber[3033] = 2'd0;
    assign memnumber[3034] = 2'd0;
    assign memnumber[3035] = 2'd0;
    assign memnumber[3036] = 2'd0;
    assign memnumber[3037] = 2'd0;
    assign memnumber[3038] = 2'd2;
    assign memnumber[3039] = 2'd2;
    assign memnumber[3040] = 2'd1;
    assign memnumber[3041] = 2'd0;
    assign memnumber[3042] = 2'd0;
    assign memnumber[3043] = 2'd0;
    assign memnumber[3044] = 2'd0;
    assign memnumber[3045] = 2'd0;
    assign memnumber[3046] = 2'd0;
    assign memnumber[3047] = 2'd0;
    assign memnumber[3048] = 2'd0;
    assign memnumber[3049] = 2'd0;
    assign memnumber[3050] = 2'd2;
    assign memnumber[3051] = 2'd2;
    assign memnumber[3052] = 2'd1;
    assign memnumber[3053] = 2'd1;
    assign memnumber[3054] = 2'd0;
    assign memnumber[3055] = 2'd0;
    assign memnumber[3056] = 2'd0;
    assign memnumber[3057] = 2'd0;
    assign memnumber[3058] = 2'd0;
    assign memnumber[3059] = 2'd0;
    assign memnumber[3060] = 2'd0;
    assign memnumber[3061] = 2'd2;
    assign memnumber[3062] = 2'd2;
    assign memnumber[3063] = 2'd1;
    assign memnumber[3064] = 2'd0;
    assign memnumber[3065] = 2'd0;
    assign memnumber[3066] = 2'd0;
    assign memnumber[3067] = 2'd0;
    assign memnumber[3068] = 2'd0;
    assign memnumber[3069] = 2'd0;
    assign memnumber[3070] = 2'd0;
    assign memnumber[3071] = 2'd0;
    assign memnumber[3072] = 2'd0;
    assign memnumber[3073] = 2'd2;
    assign memnumber[3074] = 2'd2;
    assign memnumber[3075] = 2'd1;
    assign memnumber[3076] = 2'd0;
    assign memnumber[3077] = 2'd0;
    assign memnumber[3078] = 2'd0;
    assign memnumber[3079] = 2'd0;
    assign memnumber[3080] = 2'd0;
    assign memnumber[3081] = 2'd0;
    assign memnumber[3082] = 2'd0;
    assign memnumber[3083] = 2'd0;
    assign memnumber[3084] = 2'd0;
    assign memnumber[3085] = 2'd0;
    assign memnumber[3086] = 2'd2;
    assign memnumber[3087] = 2'd2;
    assign memnumber[3088] = 2'd1;
    assign memnumber[3089] = 2'd0;
    assign memnumber[3090] = 2'd0;
    assign memnumber[3091] = 2'd0;
    assign memnumber[3092] = 2'd0;
    assign memnumber[3093] = 2'd0;
    assign memnumber[3094] = 2'd0;
    assign memnumber[3095] = 2'd0;
    assign memnumber[3096] = 2'd0;
    assign memnumber[3097] = 2'd0;
    assign memnumber[3098] = 2'd0;
    assign memnumber[3099] = 2'd0;
    assign memnumber[3100] = 2'd0;
    assign memnumber[3101] = 2'd0;
    assign memnumber[3102] = 2'd2;
    assign memnumber[3103] = 2'd2;
    assign memnumber[3104] = 2'd1;
    assign memnumber[3105] = 2'd1;
    assign memnumber[3106] = 2'd0;
    assign memnumber[3107] = 2'd0;
    assign memnumber[3108] = 2'd0;
    assign memnumber[3109] = 2'd0;
    assign memnumber[3110] = 2'd0;
    assign memnumber[3111] = 2'd0;
    assign memnumber[3112] = 2'd0;
    assign memnumber[3113] = 2'd0;
    assign memnumber[3114] = 2'd2;
    assign memnumber[3115] = 2'd2;
    assign memnumber[3116] = 2'd1;
    assign memnumber[3117] = 2'd0;
    assign memnumber[3118] = 2'd0;
    assign memnumber[3119] = 2'd0;
    assign memnumber[3120] = 2'd0;
    assign memnumber[3121] = 2'd0;
    assign memnumber[3122] = 2'd0;
    assign memnumber[3123] = 2'd0;
    assign memnumber[3124] = 2'd0;
    assign memnumber[3125] = 2'd0;
    assign memnumber[3126] = 2'd0;
    assign memnumber[3127] = 2'd0;
    assign memnumber[3128] = 2'd2;
    assign memnumber[3129] = 2'd2;
    assign memnumber[3130] = 2'd1;
    assign memnumber[3131] = 2'd0;
    assign memnumber[3132] = 2'd2;
    assign memnumber[3133] = 2'd2;
    assign memnumber[3134] = 2'd2;
    assign memnumber[3135] = 2'd2;
    assign memnumber[3136] = 2'd2;
    assign memnumber[3137] = 2'd2;
    assign memnumber[3138] = 2'd2;
    assign memnumber[3139] = 2'd2;
    assign memnumber[3140] = 2'd2;
    assign memnumber[3141] = 2'd2;
    assign memnumber[3142] = 2'd2;
    assign memnumber[3143] = 2'd2;
    assign memnumber[3144] = 2'd2;
    assign memnumber[3145] = 2'd2;
    assign memnumber[3146] = 2'd2;
    assign memnumber[3147] = 2'd2;
    assign memnumber[3148] = 2'd1;
    assign memnumber[3149] = 2'd0;
    assign memnumber[3150] = 2'd2;
    assign memnumber[3151] = 2'd2;
    assign memnumber[3152] = 2'd0;
    assign memnumber[3153] = 2'd0;
    assign memnumber[3154] = 2'd0;
    assign memnumber[3155] = 2'd0;
    assign memnumber[3156] = 2'd0;
    assign memnumber[3157] = 2'd0;
    assign memnumber[3158] = 2'd0;
    assign memnumber[3159] = 2'd0;
    assign memnumber[3160] = 2'd0;
    assign memnumber[3161] = 2'd0;
    assign memnumber[3162] = 2'd0;
    assign memnumber[3163] = 2'd2;
    assign memnumber[3164] = 2'd2;
    assign memnumber[3165] = 2'd1;
    assign memnumber[3166] = 2'd0;
    assign memnumber[3167] = 2'd0;
    assign memnumber[3168] = 2'd0;
    assign memnumber[3169] = 2'd2;
    assign memnumber[3170] = 2'd2;
    assign memnumber[3171] = 2'd1;
    assign memnumber[3172] = 2'd0;
    assign memnumber[3173] = 2'd0;
    assign memnumber[3174] = 2'd0;
    assign memnumber[3175] = 2'd0;
    assign memnumber[3176] = 2'd0;
    assign memnumber[3177] = 2'd0;
    assign memnumber[3178] = 2'd0;
    assign memnumber[3179] = 2'd0;
    assign memnumber[3180] = 2'd0;
    assign memnumber[3181] = 2'd2;
    assign memnumber[3182] = 2'd2;
    assign memnumber[3183] = 2'd1;
    assign memnumber[3184] = 2'd0;
    assign memnumber[3185] = 2'd0;
    assign memnumber[3186] = 2'd0;
    assign memnumber[3187] = 2'd0;
    assign memnumber[3188] = 2'd0;
    assign memnumber[3189] = 2'd0;
    assign memnumber[3190] = 2'd0;
    assign memnumber[3191] = 2'd2;
    assign memnumber[3192] = 2'd2;
    assign memnumber[3193] = 2'd1;
    assign memnumber[3194] = 2'd0;
    assign memnumber[3195] = 2'd0;
    assign memnumber[3196] = 2'd0;
    assign memnumber[3197] = 2'd0;
    assign memnumber[3198] = 2'd0;
    assign memnumber[3199] = 2'd0;
    assign memnumber[3200] = 2'd0;
    assign memnumber[3201] = 2'd0;
    assign memnumber[3202] = 2'd0;
    assign memnumber[3203] = 2'd0;
    assign memnumber[3204] = 2'd2;
    assign memnumber[3205] = 2'd2;
    assign memnumber[3206] = 2'd1;
    assign memnumber[3207] = 2'd0;
    assign memnumber[3208] = 2'd0;
    assign memnumber[3209] = 2'd0;
    assign memnumber[3210] = 2'd0;
    assign memnumber[3211] = 2'd0;
    assign memnumber[3212] = 2'd0;
    assign memnumber[3213] = 2'd0;
    assign memnumber[3214] = 2'd0;
    assign memnumber[3215] = 2'd0;
    assign memnumber[3216] = 2'd0;
    assign memnumber[3217] = 2'd0;
    assign memnumber[3218] = 2'd2;
    assign memnumber[3219] = 2'd2;
    assign memnumber[3220] = 2'd1;
    assign memnumber[3221] = 2'd0;
    assign memnumber[3222] = 2'd0;
    assign memnumber[3223] = 2'd0;
    assign memnumber[3224] = 2'd0;
    assign memnumber[3225] = 2'd0;
    assign memnumber[3226] = 2'd0;
    assign memnumber[3227] = 2'd0;
    assign memnumber[3228] = 2'd0;
    assign memnumber[3229] = 2'd2;
    assign memnumber[3230] = 2'd2;
    assign memnumber[3231] = 2'd1;
    assign memnumber[3232] = 2'd1;
    assign memnumber[3233] = 2'd0;
    assign memnumber[3234] = 2'd0;
    assign memnumber[3235] = 2'd0;
    assign memnumber[3236] = 2'd0;
    assign memnumber[3237] = 2'd0;
    assign memnumber[3238] = 2'd0;
    assign memnumber[3239] = 2'd0;
    assign memnumber[3240] = 2'd0;
    assign memnumber[3241] = 2'd2;
    assign memnumber[3242] = 2'd2;
    assign memnumber[3243] = 2'd1;
    assign memnumber[3244] = 2'd0;
    assign memnumber[3245] = 2'd0;
    assign memnumber[3246] = 2'd0;
    assign memnumber[3247] = 2'd0;
    assign memnumber[3248] = 2'd0;
    assign memnumber[3249] = 2'd0;
    assign memnumber[3250] = 2'd0;
    assign memnumber[3251] = 2'd0;
    assign memnumber[3252] = 2'd2;
    assign memnumber[3253] = 2'd2;
    assign memnumber[3254] = 2'd2;
    assign memnumber[3255] = 2'd1;
    assign memnumber[3256] = 2'd0;
    assign memnumber[3257] = 2'd0;
    assign memnumber[3258] = 2'd0;
    assign memnumber[3259] = 2'd0;
    assign memnumber[3260] = 2'd0;
    assign memnumber[3261] = 2'd0;
    assign memnumber[3262] = 2'd0;
    assign memnumber[3263] = 2'd0;
    assign memnumber[3264] = 2'd0;
    assign memnumber[3265] = 2'd0;
    assign memnumber[3266] = 2'd2;
    assign memnumber[3267] = 2'd2;
    assign memnumber[3268] = 2'd1;
    assign memnumber[3269] = 2'd0;
    assign memnumber[3270] = 2'd0;
    assign memnumber[3271] = 2'd0;
    assign memnumber[3272] = 2'd0;
    assign memnumber[3273] = 2'd0;
    assign memnumber[3274] = 2'd0;
    assign memnumber[3275] = 2'd0;
    assign memnumber[3276] = 2'd0;
    assign memnumber[3277] = 2'd0;
    assign memnumber[3278] = 2'd0;
    assign memnumber[3279] = 2'd0;
    assign memnumber[3280] = 2'd0;
    assign memnumber[3281] = 2'd2;
    assign memnumber[3282] = 2'd2;
    assign memnumber[3283] = 2'd1;
    assign memnumber[3284] = 2'd1;
    assign memnumber[3285] = 2'd0;
    assign memnumber[3286] = 2'd0;
    assign memnumber[3287] = 2'd0;
    assign memnumber[3288] = 2'd0;
    assign memnumber[3289] = 2'd0;
    assign memnumber[3290] = 2'd0;
    assign memnumber[3291] = 2'd0;
    assign memnumber[3292] = 2'd0;
    assign memnumber[3293] = 2'd0;
    assign memnumber[3294] = 2'd0;
    assign memnumber[3295] = 2'd2;
    assign memnumber[3296] = 2'd2;
    assign memnumber[3297] = 2'd0;
    assign memnumber[3298] = 2'd0;
    assign memnumber[3299] = 2'd0;
    assign memnumber[3300] = 2'd0;
    assign memnumber[3301] = 2'd0;
    assign memnumber[3302] = 2'd0;
    assign memnumber[3303] = 2'd0;
    assign memnumber[3304] = 2'd0;
    assign memnumber[3305] = 2'd0;
    assign memnumber[3306] = 2'd0;
    assign memnumber[3307] = 2'd2;
    assign memnumber[3308] = 2'd2;
    assign memnumber[3309] = 2'd1;
    assign memnumber[3310] = 2'd1;
    assign memnumber[3311] = 2'd0;
    assign memnumber[3312] = 2'd0;
    assign memnumber[3313] = 2'd1;
    assign memnumber[3314] = 2'd1;
    assign memnumber[3315] = 2'd1;
    assign memnumber[3316] = 2'd1;
    assign memnumber[3317] = 2'd1;
    assign memnumber[3318] = 2'd1;
    assign memnumber[3319] = 2'd1;
    assign memnumber[3320] = 2'd1;
    assign memnumber[3321] = 2'd1;
    assign memnumber[3322] = 2'd1;
    assign memnumber[3323] = 2'd2;
    assign memnumber[3324] = 2'd2;
    assign memnumber[3325] = 2'd1;
    assign memnumber[3326] = 2'd1;
    assign memnumber[3327] = 2'd1;
    assign memnumber[3328] = 2'd1;
    assign memnumber[3329] = 2'd0;
    assign memnumber[3330] = 2'd2;
    assign memnumber[3331] = 2'd2;
    assign memnumber[3332] = 2'd2;
    assign memnumber[3333] = 2'd0;
    assign memnumber[3334] = 2'd0;
    assign memnumber[3335] = 2'd0;
    assign memnumber[3336] = 2'd0;
    assign memnumber[3337] = 2'd0;
    assign memnumber[3338] = 2'd0;
    assign memnumber[3339] = 2'd0;
    assign memnumber[3340] = 2'd0;
    assign memnumber[3341] = 2'd0;
    assign memnumber[3342] = 2'd2;
    assign memnumber[3343] = 2'd2;
    assign memnumber[3344] = 2'd1;
    assign memnumber[3345] = 2'd1;
    assign memnumber[3346] = 2'd0;
    assign memnumber[3347] = 2'd0;
    assign memnumber[3348] = 2'd0;
    assign memnumber[3349] = 2'd2;
    assign memnumber[3350] = 2'd2;
    assign memnumber[3351] = 2'd2;
    assign memnumber[3352] = 2'd0;
    assign memnumber[3353] = 2'd0;
    assign memnumber[3354] = 2'd0;
    assign memnumber[3355] = 2'd0;
    assign memnumber[3356] = 2'd0;
    assign memnumber[3357] = 2'd0;
    assign memnumber[3358] = 2'd0;
    assign memnumber[3359] = 2'd0;
    assign memnumber[3360] = 2'd0;
    assign memnumber[3361] = 2'd2;
    assign memnumber[3362] = 2'd2;
    assign memnumber[3363] = 2'd1;
    assign memnumber[3364] = 2'd0;
    assign memnumber[3365] = 2'd0;
    assign memnumber[3366] = 2'd0;
    assign memnumber[3367] = 2'd0;
    assign memnumber[3368] = 2'd0;
    assign memnumber[3369] = 2'd0;
    assign memnumber[3370] = 2'd2;
    assign memnumber[3371] = 2'd2;
    assign memnumber[3372] = 2'd1;
    assign memnumber[3373] = 2'd1;
    assign memnumber[3374] = 2'd0;
    assign memnumber[3375] = 2'd0;
    assign memnumber[3376] = 2'd0;
    assign memnumber[3377] = 2'd0;
    assign memnumber[3378] = 2'd0;
    assign memnumber[3379] = 2'd0;
    assign memnumber[3380] = 2'd0;
    assign memnumber[3381] = 2'd0;
    assign memnumber[3382] = 2'd0;
    assign memnumber[3383] = 2'd0;
    assign memnumber[3384] = 2'd2;
    assign memnumber[3385] = 2'd2;
    assign memnumber[3386] = 2'd2;
    assign memnumber[3387] = 2'd0;
    assign memnumber[3388] = 2'd0;
    assign memnumber[3389] = 2'd0;
    assign memnumber[3390] = 2'd0;
    assign memnumber[3391] = 2'd0;
    assign memnumber[3392] = 2'd0;
    assign memnumber[3393] = 2'd0;
    assign memnumber[3394] = 2'd0;
    assign memnumber[3395] = 2'd0;
    assign memnumber[3396] = 2'd0;
    assign memnumber[3397] = 2'd2;
    assign memnumber[3398] = 2'd2;
    assign memnumber[3399] = 2'd1;
    assign memnumber[3400] = 2'd1;
    assign memnumber[3401] = 2'd0;
    assign memnumber[3402] = 2'd0;
    assign memnumber[3403] = 2'd0;
    assign memnumber[3404] = 2'd0;
    assign memnumber[3405] = 2'd0;
    assign memnumber[3406] = 2'd0;
    assign memnumber[3407] = 2'd0;
    assign memnumber[3408] = 2'd2;
    assign memnumber[3409] = 2'd2;
    assign memnumber[3410] = 2'd1;
    assign memnumber[3411] = 2'd1;
    assign memnumber[3412] = 2'd0;
    assign memnumber[3413] = 2'd0;
    assign memnumber[3414] = 2'd0;
    assign memnumber[3415] = 2'd0;
    assign memnumber[3416] = 2'd0;
    assign memnumber[3417] = 2'd0;
    assign memnumber[3418] = 2'd0;
    assign memnumber[3419] = 2'd0;
    assign memnumber[3420] = 2'd0;
    assign memnumber[3421] = 2'd0;
    assign memnumber[3422] = 2'd2;
    assign memnumber[3423] = 2'd2;
    assign memnumber[3424] = 2'd0;
    assign memnumber[3425] = 2'd0;
    assign memnumber[3426] = 2'd0;
    assign memnumber[3427] = 2'd0;
    assign memnumber[3428] = 2'd0;
    assign memnumber[3429] = 2'd0;
    assign memnumber[3430] = 2'd0;
    assign memnumber[3431] = 2'd0;
    assign memnumber[3432] = 2'd2;
    assign memnumber[3433] = 2'd2;
    assign memnumber[3434] = 2'd1;
    assign memnumber[3435] = 2'd1;
    assign memnumber[3436] = 2'd0;
    assign memnumber[3437] = 2'd0;
    assign memnumber[3438] = 2'd0;
    assign memnumber[3439] = 2'd0;
    assign memnumber[3440] = 2'd0;
    assign memnumber[3441] = 2'd0;
    assign memnumber[3442] = 2'd0;
    assign memnumber[3443] = 2'd0;
    assign memnumber[3444] = 2'd0;
    assign memnumber[3445] = 2'd0;
    assign memnumber[3446] = 2'd2;
    assign memnumber[3447] = 2'd2;
    assign memnumber[3448] = 2'd1;
    assign memnumber[3449] = 2'd0;
    assign memnumber[3450] = 2'd0;
    assign memnumber[3451] = 2'd0;
    assign memnumber[3452] = 2'd0;
    assign memnumber[3453] = 2'd0;
    assign memnumber[3454] = 2'd0;
    assign memnumber[3455] = 2'd0;
    assign memnumber[3456] = 2'd0;
    assign memnumber[3457] = 2'd0;
    assign memnumber[3458] = 2'd0;
    assign memnumber[3459] = 2'd0;
    assign memnumber[3460] = 2'd2;
    assign memnumber[3461] = 2'd2;
    assign memnumber[3462] = 2'd1;
    assign memnumber[3463] = 2'd1;
    assign memnumber[3464] = 2'd0;
    assign memnumber[3465] = 2'd0;
    assign memnumber[3466] = 2'd0;
    assign memnumber[3467] = 2'd0;
    assign memnumber[3468] = 2'd0;
    assign memnumber[3469] = 2'd0;
    assign memnumber[3470] = 2'd0;
    assign memnumber[3471] = 2'd0;
    assign memnumber[3472] = 2'd0;
    assign memnumber[3473] = 2'd0;
    assign memnumber[3474] = 2'd0;
    assign memnumber[3475] = 2'd2;
    assign memnumber[3476] = 2'd2;
    assign memnumber[3477] = 2'd2;
    assign memnumber[3478] = 2'd0;
    assign memnumber[3479] = 2'd0;
    assign memnumber[3480] = 2'd0;
    assign memnumber[3481] = 2'd0;
    assign memnumber[3482] = 2'd0;
    assign memnumber[3483] = 2'd0;
    assign memnumber[3484] = 2'd0;
    assign memnumber[3485] = 2'd0;
    assign memnumber[3486] = 2'd2;
    assign memnumber[3487] = 2'd2;
    assign memnumber[3488] = 2'd2;
    assign memnumber[3489] = 2'd1;
    assign memnumber[3490] = 2'd0;
    assign memnumber[3491] = 2'd0;
    assign memnumber[3492] = 2'd0;
    assign memnumber[3493] = 2'd0;
    assign memnumber[3494] = 2'd0;
    assign memnumber[3495] = 2'd0;
    assign memnumber[3496] = 2'd0;
    assign memnumber[3497] = 2'd0;
    assign memnumber[3498] = 2'd0;
    assign memnumber[3499] = 2'd0;
    assign memnumber[3500] = 2'd0;
    assign memnumber[3501] = 2'd0;
    assign memnumber[3502] = 2'd0;
    assign memnumber[3503] = 2'd2;
    assign memnumber[3504] = 2'd2;
    assign memnumber[3505] = 2'd1;
    assign memnumber[3506] = 2'd0;
    assign memnumber[3507] = 2'd0;
    assign memnumber[3508] = 2'd0;
    assign memnumber[3509] = 2'd0;
    assign memnumber[3510] = 2'd0;
    assign memnumber[3511] = 2'd2;
    assign memnumber[3512] = 2'd2;
    assign memnumber[3513] = 2'd1;
    assign memnumber[3514] = 2'd0;
    assign memnumber[3515] = 2'd0;
    assign memnumber[3516] = 2'd0;
    assign memnumber[3517] = 2'd0;
    assign memnumber[3518] = 2'd0;
    assign memnumber[3519] = 2'd0;
    assign memnumber[3520] = 2'd0;
    assign memnumber[3521] = 2'd2;
    assign memnumber[3522] = 2'd2;
    assign memnumber[3523] = 2'd2;
    assign memnumber[3524] = 2'd1;
    assign memnumber[3525] = 2'd0;
    assign memnumber[3526] = 2'd0;
    assign memnumber[3527] = 2'd0;
    assign memnumber[3528] = 2'd0;
    assign memnumber[3529] = 2'd0;
    assign memnumber[3530] = 2'd2;
    assign memnumber[3531] = 2'd2;
    assign memnumber[3532] = 2'd1;
    assign memnumber[3533] = 2'd0;
    assign memnumber[3534] = 2'd0;
    assign memnumber[3535] = 2'd0;
    assign memnumber[3536] = 2'd0;
    assign memnumber[3537] = 2'd0;
    assign memnumber[3538] = 2'd0;
    assign memnumber[3539] = 2'd0;
    assign memnumber[3540] = 2'd2;
    assign memnumber[3541] = 2'd2;
    assign memnumber[3542] = 2'd1;
    assign memnumber[3543] = 2'd1;
    assign memnumber[3544] = 2'd0;
    assign memnumber[3545] = 2'd0;
    assign memnumber[3546] = 2'd0;
    assign memnumber[3547] = 2'd0;
    assign memnumber[3548] = 2'd0;
    assign memnumber[3549] = 2'd0;
    assign memnumber[3550] = 2'd2;
    assign memnumber[3551] = 2'd2;
    assign memnumber[3552] = 2'd1;
    assign memnumber[3553] = 2'd0;
    assign memnumber[3554] = 2'd0;
    assign memnumber[3555] = 2'd0;
    assign memnumber[3556] = 2'd0;
    assign memnumber[3557] = 2'd0;
    assign memnumber[3558] = 2'd0;
    assign memnumber[3559] = 2'd0;
    assign memnumber[3560] = 2'd0;
    assign memnumber[3561] = 2'd0;
    assign memnumber[3562] = 2'd0;
    assign memnumber[3563] = 2'd0;
    assign memnumber[3564] = 2'd0;
    assign memnumber[3565] = 2'd2;
    assign memnumber[3566] = 2'd2;
    assign memnumber[3567] = 2'd1;
    assign memnumber[3568] = 2'd0;
    assign memnumber[3569] = 2'd0;
    assign memnumber[3570] = 2'd0;
    assign memnumber[3571] = 2'd0;
    assign memnumber[3572] = 2'd0;
    assign memnumber[3573] = 2'd0;
    assign memnumber[3574] = 2'd0;
    assign memnumber[3575] = 2'd0;
    assign memnumber[3576] = 2'd2;
    assign memnumber[3577] = 2'd2;
    assign memnumber[3578] = 2'd2;
    assign memnumber[3579] = 2'd1;
    assign memnumber[3580] = 2'd0;
    assign memnumber[3581] = 2'd0;
    assign memnumber[3582] = 2'd0;
    assign memnumber[3583] = 2'd0;
    assign memnumber[3584] = 2'd0;
    assign memnumber[3585] = 2'd0;
    assign memnumber[3586] = 2'd0;
    assign memnumber[3587] = 2'd2;
    assign memnumber[3588] = 2'd2;
    assign memnumber[3589] = 2'd2;
    assign memnumber[3590] = 2'd1;
    assign memnumber[3591] = 2'd0;
    assign memnumber[3592] = 2'd0;
    assign memnumber[3593] = 2'd0;
    assign memnumber[3594] = 2'd0;
    assign memnumber[3595] = 2'd0;
    assign memnumber[3596] = 2'd0;
    assign memnumber[3597] = 2'd0;
    assign memnumber[3598] = 2'd0;
    assign memnumber[3599] = 2'd0;
    assign memnumber[3600] = 2'd0;
    assign memnumber[3601] = 2'd0;
    assign memnumber[3602] = 2'd2;
    assign memnumber[3603] = 2'd2;
    assign memnumber[3604] = 2'd2;
    assign memnumber[3605] = 2'd2;
    assign memnumber[3606] = 2'd0;
    assign memnumber[3607] = 2'd0;
    assign memnumber[3608] = 2'd0;
    assign memnumber[3609] = 2'd0;
    assign memnumber[3610] = 2'd2;
    assign memnumber[3611] = 2'd2;
    assign memnumber[3612] = 2'd2;
    assign memnumber[3613] = 2'd1;
    assign memnumber[3614] = 2'd1;
    assign memnumber[3615] = 2'd0;
    assign memnumber[3616] = 2'd0;
    assign memnumber[3617] = 2'd0;
    assign memnumber[3618] = 2'd0;
    assign memnumber[3619] = 2'd0;
    assign memnumber[3620] = 2'd0;
    assign memnumber[3621] = 2'd0;
    assign memnumber[3622] = 2'd0;
    assign memnumber[3623] = 2'd0;
    assign memnumber[3624] = 2'd0;
    assign memnumber[3625] = 2'd0;
    assign memnumber[3626] = 2'd2;
    assign memnumber[3627] = 2'd2;
    assign memnumber[3628] = 2'd1;
    assign memnumber[3629] = 2'd0;
    assign memnumber[3630] = 2'd0;
    assign memnumber[3631] = 2'd0;
    assign memnumber[3632] = 2'd0;
    assign memnumber[3633] = 2'd0;
    assign memnumber[3634] = 2'd0;
    assign memnumber[3635] = 2'd0;
    assign memnumber[3636] = 2'd0;
    assign memnumber[3637] = 2'd0;
    assign memnumber[3638] = 2'd0;
    assign memnumber[3639] = 2'd2;
    assign memnumber[3640] = 2'd2;
    assign memnumber[3641] = 2'd1;
    assign memnumber[3642] = 2'd1;
    assign memnumber[3643] = 2'd0;
    assign memnumber[3644] = 2'd0;
    assign memnumber[3645] = 2'd0;
    assign memnumber[3646] = 2'd0;
    assign memnumber[3647] = 2'd0;
    assign memnumber[3648] = 2'd0;
    assign memnumber[3649] = 2'd0;
    assign memnumber[3650] = 2'd0;
    assign memnumber[3651] = 2'd0;
    assign memnumber[3652] = 2'd0;
    assign memnumber[3653] = 2'd0;
    assign memnumber[3654] = 2'd0;
    assign memnumber[3655] = 2'd0;
    assign memnumber[3656] = 2'd2;
    assign memnumber[3657] = 2'd2;
    assign memnumber[3658] = 2'd2;
    assign memnumber[3659] = 2'd0;
    assign memnumber[3660] = 2'd0;
    assign memnumber[3661] = 2'd0;
    assign memnumber[3662] = 2'd0;
    assign memnumber[3663] = 2'd0;
    assign memnumber[3664] = 2'd0;
    assign memnumber[3665] = 2'd2;
    assign memnumber[3666] = 2'd2;
    assign memnumber[3667] = 2'd2;
    assign memnumber[3668] = 2'd1;
    assign memnumber[3669] = 2'd1;
    assign memnumber[3670] = 2'd0;
    assign memnumber[3671] = 2'd0;
    assign memnumber[3672] = 2'd0;
    assign memnumber[3673] = 2'd0;
    assign memnumber[3674] = 2'd0;
    assign memnumber[3675] = 2'd0;
    assign memnumber[3676] = 2'd0;
    assign memnumber[3677] = 2'd0;
    assign memnumber[3678] = 2'd0;
    assign memnumber[3679] = 2'd0;
    assign memnumber[3680] = 2'd0;
    assign memnumber[3681] = 2'd0;
    assign memnumber[3682] = 2'd0;
    assign memnumber[3683] = 2'd2;
    assign memnumber[3684] = 2'd2;
    assign memnumber[3685] = 2'd1;
    assign memnumber[3686] = 2'd0;
    assign memnumber[3687] = 2'd0;
    assign memnumber[3688] = 2'd0;
    assign memnumber[3689] = 2'd0;
    assign memnumber[3690] = 2'd0;
    assign memnumber[3691] = 2'd2;
    assign memnumber[3692] = 2'd2;
    assign memnumber[3693] = 2'd2;
    assign memnumber[3694] = 2'd2;
    assign memnumber[3695] = 2'd0;
    assign memnumber[3696] = 2'd0;
    assign memnumber[3697] = 2'd0;
    assign memnumber[3698] = 2'd0;
    assign memnumber[3699] = 2'd0;
    assign memnumber[3700] = 2'd2;
    assign memnumber[3701] = 2'd2;
    assign memnumber[3702] = 2'd2;
    assign memnumber[3703] = 2'd1;
    assign memnumber[3704] = 2'd1;
    assign memnumber[3705] = 2'd0;
    assign memnumber[3706] = 2'd0;
    assign memnumber[3707] = 2'd0;
    assign memnumber[3708] = 2'd0;
    assign memnumber[3709] = 2'd0;
    assign memnumber[3710] = 2'd2;
    assign memnumber[3711] = 2'd2;
    assign memnumber[3712] = 2'd2;
    assign memnumber[3713] = 2'd2;
    assign memnumber[3714] = 2'd0;
    assign memnumber[3715] = 2'd0;
    assign memnumber[3716] = 2'd0;
    assign memnumber[3717] = 2'd0;
    assign memnumber[3718] = 2'd2;
    assign memnumber[3719] = 2'd2;
    assign memnumber[3720] = 2'd2;
    assign memnumber[3721] = 2'd2;
    assign memnumber[3722] = 2'd1;
    assign memnumber[3723] = 2'd0;
    assign memnumber[3724] = 2'd0;
    assign memnumber[3725] = 2'd0;
    assign memnumber[3726] = 2'd0;
    assign memnumber[3727] = 2'd0;
    assign memnumber[3728] = 2'd0;
    assign memnumber[3729] = 2'd2;
    assign memnumber[3730] = 2'd2;
    assign memnumber[3731] = 2'd1;
    assign memnumber[3732] = 2'd1;
    assign memnumber[3733] = 2'd0;
    assign memnumber[3734] = 2'd0;
    assign memnumber[3735] = 2'd0;
    assign memnumber[3736] = 2'd0;
    assign memnumber[3737] = 2'd0;
    assign memnumber[3738] = 2'd0;
    assign memnumber[3739] = 2'd0;
    assign memnumber[3740] = 2'd0;
    assign memnumber[3741] = 2'd0;
    assign memnumber[3742] = 2'd0;
    assign memnumber[3743] = 2'd0;
    assign memnumber[3744] = 2'd0;
    assign memnumber[3745] = 2'd0;
    assign memnumber[3746] = 2'd2;
    assign memnumber[3747] = 2'd2;
    assign memnumber[3748] = 2'd2;
    assign memnumber[3749] = 2'd0;
    assign memnumber[3750] = 2'd0;
    assign memnumber[3751] = 2'd0;
    assign memnumber[3752] = 2'd0;
    assign memnumber[3753] = 2'd0;
    assign memnumber[3754] = 2'd0;
    assign memnumber[3755] = 2'd2;
    assign memnumber[3756] = 2'd2;
    assign memnumber[3757] = 2'd2;
    assign memnumber[3758] = 2'd1;
    assign memnumber[3759] = 2'd1;
    assign memnumber[3760] = 2'd0;
    assign memnumber[3761] = 2'd0;
    assign memnumber[3762] = 2'd0;
    assign memnumber[3763] = 2'd0;
    assign memnumber[3764] = 2'd0;
    assign memnumber[3765] = 2'd0;
    assign memnumber[3766] = 2'd0;
    assign memnumber[3767] = 2'd2;
    assign memnumber[3768] = 2'd2;
    assign memnumber[3769] = 2'd1;
    assign memnumber[3770] = 2'd1;
    assign memnumber[3771] = 2'd0;
    assign memnumber[3772] = 2'd0;
    assign memnumber[3773] = 2'd0;
    assign memnumber[3774] = 2'd0;
    assign memnumber[3775] = 2'd0;
    assign memnumber[3776] = 2'd0;
    assign memnumber[3777] = 2'd0;
    assign memnumber[3778] = 2'd0;
    assign memnumber[3779] = 2'd0;
    assign memnumber[3780] = 2'd0;
    assign memnumber[3781] = 2'd0;
    assign memnumber[3782] = 2'd0;
    assign memnumber[3783] = 2'd2;
    assign memnumber[3784] = 2'd2;
    assign memnumber[3785] = 2'd2;
    assign memnumber[3786] = 2'd2;
    assign memnumber[3787] = 2'd2;
    assign memnumber[3788] = 2'd2;
    assign memnumber[3789] = 2'd2;
    assign memnumber[3790] = 2'd2;
    assign memnumber[3791] = 2'd2;
    assign memnumber[3792] = 2'd1;
    assign memnumber[3793] = 2'd1;
    assign memnumber[3794] = 2'd0;
    assign memnumber[3795] = 2'd0;
    assign memnumber[3796] = 2'd0;
    assign memnumber[3797] = 2'd0;
    assign memnumber[3798] = 2'd0;
    assign memnumber[3799] = 2'd0;
    assign memnumber[3800] = 2'd0;
    assign memnumber[3801] = 2'd0;
    assign memnumber[3802] = 2'd0;
    assign memnumber[3803] = 2'd0;
    assign memnumber[3804] = 2'd0;
    assign memnumber[3805] = 2'd0;
    assign memnumber[3806] = 2'd2;
    assign memnumber[3807] = 2'd2;
    assign memnumber[3808] = 2'd1;
    assign memnumber[3809] = 2'd0;
    assign memnumber[3810] = 2'd0;
    assign memnumber[3811] = 2'd0;
    assign memnumber[3812] = 2'd0;
    assign memnumber[3813] = 2'd0;
    assign memnumber[3814] = 2'd0;
    assign memnumber[3815] = 2'd0;
    assign memnumber[3816] = 2'd0;
    assign memnumber[3817] = 2'd0;
    assign memnumber[3818] = 2'd2;
    assign memnumber[3819] = 2'd2;
    assign memnumber[3820] = 2'd2;
    assign memnumber[3821] = 2'd2;
    assign memnumber[3822] = 2'd2;
    assign memnumber[3823] = 2'd2;
    assign memnumber[3824] = 2'd2;
    assign memnumber[3825] = 2'd2;
    assign memnumber[3826] = 2'd2;
    assign memnumber[3827] = 2'd2;
    assign memnumber[3828] = 2'd2;
    assign memnumber[3829] = 2'd2;
    assign memnumber[3830] = 2'd2;
    assign memnumber[3831] = 2'd2;
    assign memnumber[3832] = 2'd0;
    assign memnumber[3833] = 2'd0;
    assign memnumber[3834] = 2'd0;
    assign memnumber[3835] = 2'd0;
    assign memnumber[3836] = 2'd0;
    assign memnumber[3837] = 2'd2;
    assign memnumber[3838] = 2'd2;
    assign memnumber[3839] = 2'd2;
    assign memnumber[3840] = 2'd2;
    assign memnumber[3841] = 2'd2;
    assign memnumber[3842] = 2'd2;
    assign memnumber[3843] = 2'd2;
    assign memnumber[3844] = 2'd2;
    assign memnumber[3845] = 2'd2;
    assign memnumber[3846] = 2'd2;
    assign memnumber[3847] = 2'd1;
    assign memnumber[3848] = 2'd1;
    assign memnumber[3849] = 2'd0;
    assign memnumber[3850] = 2'd0;
    assign memnumber[3851] = 2'd0;
    assign memnumber[3852] = 2'd0;
    assign memnumber[3853] = 2'd0;
    assign memnumber[3854] = 2'd0;
    assign memnumber[3855] = 2'd0;
    assign memnumber[3856] = 2'd0;
    assign memnumber[3857] = 2'd0;
    assign memnumber[3858] = 2'd0;
    assign memnumber[3859] = 2'd0;
    assign memnumber[3860] = 2'd0;
    assign memnumber[3861] = 2'd0;
    assign memnumber[3862] = 2'd0;
    assign memnumber[3863] = 2'd2;
    assign memnumber[3864] = 2'd2;
    assign memnumber[3865] = 2'd1;
    assign memnumber[3866] = 2'd0;
    assign memnumber[3867] = 2'd0;
    assign memnumber[3868] = 2'd0;
    assign memnumber[3869] = 2'd0;
    assign memnumber[3870] = 2'd0;
    assign memnumber[3871] = 2'd0;
    assign memnumber[3872] = 2'd1;
    assign memnumber[3873] = 2'd2;
    assign memnumber[3874] = 2'd2;
    assign memnumber[3875] = 2'd2;
    assign memnumber[3876] = 2'd2;
    assign memnumber[3877] = 2'd2;
    assign memnumber[3878] = 2'd2;
    assign memnumber[3879] = 2'd2;
    assign memnumber[3880] = 2'd2;
    assign memnumber[3881] = 2'd2;
    assign memnumber[3882] = 2'd1;
    assign memnumber[3883] = 2'd1;
    assign memnumber[3884] = 2'd0;
    assign memnumber[3885] = 2'd0;
    assign memnumber[3886] = 2'd0;
    assign memnumber[3887] = 2'd0;
    assign memnumber[3888] = 2'd0;
    assign memnumber[3889] = 2'd0;
    assign memnumber[3890] = 2'd0;
    assign memnumber[3891] = 2'd2;
    assign memnumber[3892] = 2'd2;
    assign memnumber[3893] = 2'd2;
    assign memnumber[3894] = 2'd2;
    assign memnumber[3895] = 2'd2;
    assign memnumber[3896] = 2'd2;
    assign memnumber[3897] = 2'd2;
    assign memnumber[3898] = 2'd2;
    assign memnumber[3899] = 2'd2;
    assign memnumber[3900] = 2'd1;
    assign memnumber[3901] = 2'd1;
    assign memnumber[3902] = 2'd1;
    assign memnumber[3903] = 2'd0;
    assign memnumber[3904] = 2'd0;
    assign memnumber[3905] = 2'd0;
    assign memnumber[3906] = 2'd0;
    assign memnumber[3907] = 2'd0;
    assign memnumber[3908] = 2'd0;
    assign memnumber[3909] = 2'd2;
    assign memnumber[3910] = 2'd2;
    assign memnumber[3911] = 2'd1;
    assign memnumber[3912] = 2'd0;
    assign memnumber[3913] = 2'd0;
    assign memnumber[3914] = 2'd0;
    assign memnumber[3915] = 2'd0;
    assign memnumber[3916] = 2'd0;
    assign memnumber[3917] = 2'd0;
    assign memnumber[3918] = 2'd0;
    assign memnumber[3919] = 2'd0;
    assign memnumber[3920] = 2'd0;
    assign memnumber[3921] = 2'd0;
    assign memnumber[3922] = 2'd0;
    assign memnumber[3923] = 2'd0;
    assign memnumber[3924] = 2'd0;
    assign memnumber[3925] = 2'd0;
    assign memnumber[3926] = 2'd0;
    assign memnumber[3927] = 2'd2;
    assign memnumber[3928] = 2'd2;
    assign memnumber[3929] = 2'd2;
    assign memnumber[3930] = 2'd2;
    assign memnumber[3931] = 2'd2;
    assign memnumber[3932] = 2'd2;
    assign memnumber[3933] = 2'd2;
    assign memnumber[3934] = 2'd2;
    assign memnumber[3935] = 2'd2;
    assign memnumber[3936] = 2'd2;
    assign memnumber[3937] = 2'd1;
    assign memnumber[3938] = 2'd1;
    assign memnumber[3939] = 2'd0;
    assign memnumber[3940] = 2'd0;
    assign memnumber[3941] = 2'd0;
    assign memnumber[3942] = 2'd0;
    assign memnumber[3943] = 2'd0;
    assign memnumber[3944] = 2'd0;
    assign memnumber[3945] = 2'd0;
    assign memnumber[3946] = 2'd2;
    assign memnumber[3947] = 2'd2;
    assign memnumber[3948] = 2'd1;
    assign memnumber[3949] = 2'd1;
    assign memnumber[3950] = 2'd0;
    assign memnumber[3951] = 2'd0;
    assign memnumber[3952] = 2'd0;
    assign memnumber[3953] = 2'd0;
    assign memnumber[3954] = 2'd0;
    assign memnumber[3955] = 2'd0;
    assign memnumber[3956] = 2'd0;
    assign memnumber[3957] = 2'd0;
    assign memnumber[3958] = 2'd0;
    assign memnumber[3959] = 2'd0;
    assign memnumber[3960] = 2'd0;
    assign memnumber[3961] = 2'd0;
    assign memnumber[3962] = 2'd0;
    assign memnumber[3963] = 2'd0;
    assign memnumber[3964] = 2'd1;
    assign memnumber[3965] = 2'd2;
    assign memnumber[3966] = 2'd2;
    assign memnumber[3967] = 2'd2;
    assign memnumber[3968] = 2'd2;
    assign memnumber[3969] = 2'd2;
    assign memnumber[3970] = 2'd2;
    assign memnumber[3971] = 2'd1;
    assign memnumber[3972] = 2'd1;
    assign memnumber[3973] = 2'd0;
    assign memnumber[3974] = 2'd0;
    assign memnumber[3975] = 2'd0;
    assign memnumber[3976] = 2'd0;
    assign memnumber[3977] = 2'd0;
    assign memnumber[3978] = 2'd0;
    assign memnumber[3979] = 2'd0;
    assign memnumber[3980] = 2'd0;
    assign memnumber[3981] = 2'd0;
    assign memnumber[3982] = 2'd0;
    assign memnumber[3983] = 2'd0;
    assign memnumber[3984] = 2'd0;
    assign memnumber[3985] = 2'd0;
    assign memnumber[3986] = 2'd2;
    assign memnumber[3987] = 2'd2;
    assign memnumber[3988] = 2'd1;
    assign memnumber[3989] = 2'd0;
    assign memnumber[3990] = 2'd0;
    assign memnumber[3991] = 2'd0;
    assign memnumber[3992] = 2'd0;
    assign memnumber[3993] = 2'd0;
    assign memnumber[3994] = 2'd0;
    assign memnumber[3995] = 2'd0;
    assign memnumber[3996] = 2'd0;
    assign memnumber[3997] = 2'd2;
    assign memnumber[3998] = 2'd2;
    assign memnumber[3999] = 2'd2;
    assign memnumber[4000] = 2'd2;
    assign memnumber[4001] = 2'd2;
    assign memnumber[4002] = 2'd2;
    assign memnumber[4003] = 2'd2;
    assign memnumber[4004] = 2'd2;
    assign memnumber[4005] = 2'd2;
    assign memnumber[4006] = 2'd2;
    assign memnumber[4007] = 2'd2;
    assign memnumber[4008] = 2'd2;
    assign memnumber[4009] = 2'd2;
    assign memnumber[4010] = 2'd2;
    assign memnumber[4011] = 2'd2;
    assign memnumber[4012] = 2'd1;
    assign memnumber[4013] = 2'd0;
    assign memnumber[4014] = 2'd0;
    assign memnumber[4015] = 2'd0;
    assign memnumber[4016] = 2'd0;
    assign memnumber[4017] = 2'd0;
    assign memnumber[4018] = 2'd1;
    assign memnumber[4019] = 2'd2;
    assign memnumber[4020] = 2'd2;
    assign memnumber[4021] = 2'd2;
    assign memnumber[4022] = 2'd2;
    assign memnumber[4023] = 2'd2;
    assign memnumber[4024] = 2'd2;
    assign memnumber[4025] = 2'd1;
    assign memnumber[4026] = 2'd1;
    assign memnumber[4027] = 2'd1;
    assign memnumber[4028] = 2'd0;
    assign memnumber[4029] = 2'd0;
    assign memnumber[4030] = 2'd0;
    assign memnumber[4031] = 2'd0;
    assign memnumber[4032] = 2'd0;
    assign memnumber[4033] = 2'd0;
    assign memnumber[4034] = 2'd0;
    assign memnumber[4035] = 2'd0;
    assign memnumber[4036] = 2'd0;
    assign memnumber[4037] = 2'd0;
    assign memnumber[4038] = 2'd0;
    assign memnumber[4039] = 2'd0;
    assign memnumber[4040] = 2'd0;
    assign memnumber[4041] = 2'd0;
    assign memnumber[4042] = 2'd0;
    assign memnumber[4043] = 2'd2;
    assign memnumber[4044] = 2'd2;
    assign memnumber[4045] = 2'd1;
    assign memnumber[4046] = 2'd0;
    assign memnumber[4047] = 2'd0;
    assign memnumber[4048] = 2'd0;
    assign memnumber[4049] = 2'd0;
    assign memnumber[4050] = 2'd0;
    assign memnumber[4051] = 2'd0;
    assign memnumber[4052] = 2'd0;
    assign memnumber[4053] = 2'd0;
    assign memnumber[4054] = 2'd2;
    assign memnumber[4055] = 2'd2;
    assign memnumber[4056] = 2'd2;
    assign memnumber[4057] = 2'd2;
    assign memnumber[4058] = 2'd2;
    assign memnumber[4059] = 2'd2;
    assign memnumber[4060] = 2'd1;
    assign memnumber[4061] = 2'd1;
    assign memnumber[4062] = 2'd1;
    assign memnumber[4063] = 2'd0;
    assign memnumber[4064] = 2'd0;
    assign memnumber[4065] = 2'd0;
    assign memnumber[4066] = 2'd0;
    assign memnumber[4067] = 2'd0;
    assign memnumber[4068] = 2'd0;
    assign memnumber[4069] = 2'd0;
    assign memnumber[4070] = 2'd0;
    assign memnumber[4071] = 2'd0;
    assign memnumber[4072] = 2'd1;
    assign memnumber[4073] = 2'd2;
    assign memnumber[4074] = 2'd2;
    assign memnumber[4075] = 2'd2;
    assign memnumber[4076] = 2'd2;
    assign memnumber[4077] = 2'd2;
    assign memnumber[4078] = 2'd2;
    assign memnumber[4079] = 2'd1;
    assign memnumber[4080] = 2'd1;
    assign memnumber[4081] = 2'd0;
    assign memnumber[4082] = 2'd0;
    assign memnumber[4083] = 2'd0;
    assign memnumber[4084] = 2'd0;
    assign memnumber[4085] = 2'd0;
    assign memnumber[4086] = 2'd0;
    assign memnumber[4087] = 2'd0;
    assign memnumber[4088] = 2'd2;
    assign memnumber[4089] = 2'd2;
    assign memnumber[4090] = 2'd1;
    assign memnumber[4091] = 2'd1;
    assign memnumber[4092] = 2'd0;
    assign memnumber[4093] = 2'd0;
    assign memnumber[4094] = 2'd0;
    assign memnumber[4095] = 2'd0;
    assign memnumber[4096] = 2'd0;
    assign memnumber[4097] = 2'd0;
    assign memnumber[4098] = 2'd0;
    assign memnumber[4099] = 2'd0;
    assign memnumber[4100] = 2'd0;
    assign memnumber[4101] = 2'd0;
    assign memnumber[4102] = 2'd0;
    assign memnumber[4103] = 2'd0;
    assign memnumber[4104] = 2'd0;
    assign memnumber[4105] = 2'd0;
    assign memnumber[4106] = 2'd0;
    assign memnumber[4107] = 2'd0;
    assign memnumber[4108] = 2'd1;
    assign memnumber[4109] = 2'd2;
    assign memnumber[4110] = 2'd2;
    assign memnumber[4111] = 2'd2;
    assign memnumber[4112] = 2'd2;
    assign memnumber[4113] = 2'd2;
    assign memnumber[4114] = 2'd2;
    assign memnumber[4115] = 2'd1;
    assign memnumber[4116] = 2'd1;
    assign memnumber[4117] = 2'd1;
    assign memnumber[4118] = 2'd0;
    assign memnumber[4119] = 2'd0;
    assign memnumber[4120] = 2'd0;
    assign memnumber[4121] = 2'd0;
    assign memnumber[4122] = 2'd0;
    assign memnumber[4123] = 2'd0;
    assign memnumber[4124] = 2'd0;
    assign memnumber[4125] = 2'd2;
    assign memnumber[4126] = 2'd2;
    assign memnumber[4127] = 2'd1;
    assign memnumber[4128] = 2'd1;
    assign memnumber[4129] = 2'd0;
    assign memnumber[4130] = 2'd0;
    assign memnumber[4131] = 2'd0;
    assign memnumber[4132] = 2'd0;
    assign memnumber[4133] = 2'd0;
    assign memnumber[4134] = 2'd0;
    assign memnumber[4135] = 2'd0;
    assign memnumber[4136] = 2'd0;
    assign memnumber[4137] = 2'd0;
    assign memnumber[4138] = 2'd0;
    assign memnumber[4139] = 2'd0;
    assign memnumber[4140] = 2'd0;
    assign memnumber[4141] = 2'd0;
    assign memnumber[4142] = 2'd0;
    assign memnumber[4143] = 2'd0;
    assign memnumber[4144] = 2'd0;
    assign memnumber[4145] = 2'd0;
    assign memnumber[4146] = 2'd1;
    assign memnumber[4147] = 2'd1;
    assign memnumber[4148] = 2'd1;
    assign memnumber[4149] = 2'd1;
    assign memnumber[4150] = 2'd1;
    assign memnumber[4151] = 2'd1;
    assign memnumber[4152] = 2'd0;
    assign memnumber[4153] = 2'd0;
    assign memnumber[4154] = 2'd0;
    assign memnumber[4155] = 2'd0;
    assign memnumber[4156] = 2'd0;
    assign memnumber[4157] = 2'd0;
    assign memnumber[4158] = 2'd0;
    assign memnumber[4159] = 2'd0;
    assign memnumber[4160] = 2'd0;
    assign memnumber[4161] = 2'd0;
    assign memnumber[4162] = 2'd0;
    assign memnumber[4163] = 2'd0;
    assign memnumber[4164] = 2'd0;
    assign memnumber[4165] = 2'd0;
    assign memnumber[4166] = 2'd0;
    assign memnumber[4167] = 2'd1;
    assign memnumber[4168] = 2'd1;
    assign memnumber[4169] = 2'd0;
    assign memnumber[4170] = 2'd0;
    assign memnumber[4171] = 2'd0;
    assign memnumber[4172] = 2'd0;
    assign memnumber[4173] = 2'd0;
    assign memnumber[4174] = 2'd0;
    assign memnumber[4175] = 2'd0;
    assign memnumber[4176] = 2'd0;
    assign memnumber[4177] = 2'd0;
    assign memnumber[4178] = 2'd1;
    assign memnumber[4179] = 2'd1;
    assign memnumber[4180] = 2'd1;
    assign memnumber[4181] = 2'd1;
    assign memnumber[4182] = 2'd1;
    assign memnumber[4183] = 2'd1;
    assign memnumber[4184] = 2'd1;
    assign memnumber[4185] = 2'd1;
    assign memnumber[4186] = 2'd1;
    assign memnumber[4187] = 2'd1;
    assign memnumber[4188] = 2'd1;
    assign memnumber[4189] = 2'd1;
    assign memnumber[4190] = 2'd1;
    assign memnumber[4191] = 2'd1;
    assign memnumber[4192] = 2'd1;
    assign memnumber[4193] = 2'd0;
    assign memnumber[4194] = 2'd0;
    assign memnumber[4195] = 2'd0;
    assign memnumber[4196] = 2'd0;
    assign memnumber[4197] = 2'd0;
    assign memnumber[4198] = 2'd0;
    assign memnumber[4199] = 2'd0;
    assign memnumber[4200] = 2'd1;
    assign memnumber[4201] = 2'd1;
    assign memnumber[4202] = 2'd1;
    assign memnumber[4203] = 2'd1;
    assign memnumber[4204] = 2'd1;
    assign memnumber[4205] = 2'd1;
    assign memnumber[4206] = 2'd0;
    assign memnumber[4207] = 2'd0;
    assign memnumber[4208] = 2'd0;
    assign memnumber[4209] = 2'd0;
    assign memnumber[4210] = 2'd0;
    assign memnumber[4211] = 2'd0;
    assign memnumber[4212] = 2'd0;
    assign memnumber[4213] = 2'd0;
    assign memnumber[4214] = 2'd0;
    assign memnumber[4215] = 2'd0;
    assign memnumber[4216] = 2'd0;
    assign memnumber[4217] = 2'd0;
    assign memnumber[4218] = 2'd0;
    assign memnumber[4219] = 2'd0;
    assign memnumber[4220] = 2'd0;
    assign memnumber[4221] = 2'd0;
    assign memnumber[4222] = 2'd0;
    assign memnumber[4223] = 2'd0;
    assign memnumber[4224] = 2'd1;
    assign memnumber[4225] = 2'd1;
    assign memnumber[4226] = 2'd0;
    assign memnumber[4227] = 2'd0;
    assign memnumber[4228] = 2'd0;
    assign memnumber[4229] = 2'd0;
    assign memnumber[4230] = 2'd0;
    assign memnumber[4231] = 2'd0;
    assign memnumber[4232] = 2'd0;
    assign memnumber[4233] = 2'd0;
    assign memnumber[4234] = 2'd0;
    assign memnumber[4235] = 2'd1;
    assign memnumber[4236] = 2'd1;
    assign memnumber[4237] = 2'd1;
    assign memnumber[4238] = 2'd1;
    assign memnumber[4239] = 2'd1;
    assign memnumber[4240] = 2'd1;
    assign memnumber[4241] = 2'd0;
    assign memnumber[4242] = 2'd0;
    assign memnumber[4243] = 2'd0;
    assign memnumber[4244] = 2'd0;
    assign memnumber[4245] = 2'd0;
    assign memnumber[4246] = 2'd0;
    assign memnumber[4247] = 2'd0;
    assign memnumber[4248] = 2'd0;
    assign memnumber[4249] = 2'd0;
    assign memnumber[4250] = 2'd0;
    assign memnumber[4251] = 2'd0;
    assign memnumber[4252] = 2'd0;
    assign memnumber[4253] = 2'd0;
    assign memnumber[4254] = 2'd1;
    assign memnumber[4255] = 2'd1;
    assign memnumber[4256] = 2'd1;
    assign memnumber[4257] = 2'd1;
    assign memnumber[4258] = 2'd1;
    assign memnumber[4259] = 2'd1;
    assign memnumber[4260] = 2'd0;
    assign memnumber[4261] = 2'd0;
    assign memnumber[4262] = 2'd0;
    assign memnumber[4263] = 2'd0;
    assign memnumber[4264] = 2'd0;
    assign memnumber[4265] = 2'd0;
    assign memnumber[4266] = 2'd0;
    assign memnumber[4267] = 2'd0;
    assign memnumber[4268] = 2'd0;
    assign memnumber[4269] = 2'd1;
    assign memnumber[4270] = 2'd1;
    assign memnumber[4271] = 2'd0;
    assign memnumber[4272] = 2'd0;
    assign memnumber[4273] = 2'd0;
    assign memnumber[4274] = 2'd0;
    assign memnumber[4275] = 2'd0;
    assign memnumber[4276] = 2'd0;
    assign memnumber[4277] = 2'd0;
    assign memnumber[4278] = 2'd0;
    assign memnumber[4279] = 2'd0;
    assign memnumber[4280] = 2'd0;
    assign memnumber[4281] = 2'd0;
    assign memnumber[4282] = 2'd0;
    assign memnumber[4283] = 2'd0;
    assign memnumber[4284] = 2'd0;
    assign memnumber[4285] = 2'd0;
    assign memnumber[4286] = 2'd0;
    assign memnumber[4287] = 2'd0;
    assign memnumber[4288] = 2'd0;
    assign memnumber[4289] = 2'd0;
    assign memnumber[4290] = 2'd1;
    assign memnumber[4291] = 2'd1;
    assign memnumber[4292] = 2'd1;
    assign memnumber[4293] = 2'd1;
    assign memnumber[4294] = 2'd1;
    assign memnumber[4295] = 2'd1;
    assign memnumber[4296] = 2'd0;
    assign memnumber[4297] = 2'd0;
    assign memnumber[4298] = 2'd0;
    assign memnumber[4299] = 2'd0;
    assign memnumber[4300] = 2'd0;
    assign memnumber[4301] = 2'd0;
    assign memnumber[4302] = 2'd0;
    assign memnumber[4303] = 2'd0;
    assign memnumber[4304] = 2'd0;
    assign memnumber[4305] = 2'd0;
    assign memnumber[4306] = 2'd1;
    assign memnumber[4307] = 2'd1;
    assign memnumber[4308] = 2'd0;
    assign memnumber[4309] = 2'd0;
    assign memnumber[4310] = 2'd0;
    assign memnumber[4311] = 2'd0;
    assign memnumber[4312] = 2'd0;
    assign memnumber[4313] = 2'd0;
    assign memnumber[4314] = 2'd0;
    assign memnumber[4315] = 2'd0;
    assign memnumber[4316] = 2'd0;
    assign memnumber[4317] = 2'd0;
    assign memnumber[4318] = 2'd0;
    assign memnumber[4319] = 2'd0;

endmodule
