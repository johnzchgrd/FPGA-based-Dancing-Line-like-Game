module image_rom (
    input clk,
    input valid,
    input type,
    input [1:0] song,
    input [5:0] x, y,
	output reg [11:0] dout
    );
	
	wire [2:0] memory1a [1023:0], memory1b [1023:0];
	wire [2:0] memory3a [1023:0], memory3b [1023:0];
	wire [2:0] memory4a [1023:0], memory4b [1023:0];
	wire [11:0] memcol1a [7:0], memcol1b [5:0];
	wire [11:0] memcol3a [4:0], memcol3b [7:0];
	wire [11:0] memcol4a [6:0], memcol4b [4:0];
	wire [9:0] pixel;
	wire [11:0] color1a, color1b, color3a, color3b, color4a, color4b;
	
	assign pixel = (y<<5)+x-2;
	assign color1a = (valid && song == 2'b00 && type == 0) ? memcol1a[memory1a[pixel]] : memcol1a[7];
	assign color1b = (valid && song == 2'b00 && type == 1) ? memcol1b[memory1b[pixel]] : memcol1b[5];
	assign color3a = (valid && song == 2'b10 && type == 0) ? memcol3a[memory3a[pixel]] : memcol3a[4];
	assign color3b = (valid && song == 2'b10 && type == 1) ? memcol3b[memory3b[pixel]] : memcol3b[7];
	assign color4a = (valid && song == 2'b11 && type == 0) ? memcol4a[memory4a[pixel]] : memcol4a[6];
    assign color4b = (valid && song == 2'b11 && type == 1) ? memcol4b[memory4b[pixel]] : memcol4b[4];

	always @(*) begin
	    if (~valid) begin
	       dout = 12'h000;
	    end else begin
            case (song)
                2'b00: dout = type ? color1b : color1a;
                2'b01: dout = type ? 12'hfff : 12'h000;
                2'b10: dout = type ? color3b : color3a;
                2'b11: dout = type ? color4b : color4a;
                default: dout = type ? 12'hfff : 12'h000;
            endcase
        end
    end

    assign memcol1a[0] = 12'h543;
    assign memcol1a[1] = 12'h764;
    assign memcol1a[2] = 12'h875;
    assign memcol1a[3] = 12'ha98;
    assign memcol1a[4] = 12'h997;
    assign memcol1a[5] = 12'h986;
    assign memcol1a[6] = 12'h987;
    assign memcol1a[7] = 12'h000;


    assign memcol1b[0] = 12'h998;
    assign memcol1b[1] = 12'h898;
    assign memcol1b[2] = 12'h888;
    assign memcol1b[3] = 12'h887;
    assign memcol1b[4] = 12'h999;
    assign memcol1b[5] = 12'h000;

    assign memcol3a[0] = 12'h670;
    assign memcol3a[1] = 12'h450;
    assign memcol3a[2] = 12'h990;
    assign memcol3a[3] = 12'h560;
    assign memcol3a[4] = 12'h000;

    assign memcol3b[0] = 12'hd84;
    assign memcol3b[1] = 12'hd74;
    assign memcol3b[2] = 12'hd85;
    assign memcol3b[3] = 12'hc94;
    assign memcol3b[4] = 12'hccc;
    assign memcol3b[5] = 12'haaa;
    assign memcol3b[6] = 12'hbe1;
    assign memcol3b[7] = 12'h000;

    assign memcol4a[0] = 12'h300;
    assign memcol4a[1] = 12'h401;
    assign memcol4a[2] = 12'h501;
    assign memcol4a[3] = 12'hfe0;
    assign memcol4a[4] = 12'haaa;
    assign memcol4a[5] = 12'heeb;
    assign memcol4a[6] = 12'h000;

    assign memcol4b[0] = 12'h654;
    assign memcol4b[1] = 12'h898;
    assign memcol4b[2] = 12'hcbb;
    assign memcol4b[3] = 12'haba;
    assign memcol4b[4] = 12'h000;

    assign memory1a[0   ] = 3'd0;
    assign memory1a[1   ] = 3'd0;
    assign memory1a[2   ] = 3'd0;
    assign memory1a[3   ] = 3'd0;
    assign memory1a[4   ] = 3'd0;
    assign memory1a[5   ] = 3'd1;
    assign memory1a[6   ] = 3'd1;
    assign memory1a[7   ] = 3'd0;
    assign memory1a[8   ] = 3'd0;
    assign memory1a[9   ] = 3'd0;
    assign memory1a[10  ] = 3'd0;
    assign memory1a[11  ] = 3'd0;
    assign memory1a[12  ] = 3'd0;
    assign memory1a[13  ] = 3'd1;
    assign memory1a[14  ] = 3'd0;
    assign memory1a[15  ] = 3'd0;
    assign memory1a[16  ] = 3'd0;
    assign memory1a[17  ] = 3'd0;
    assign memory1a[18  ] = 3'd0;
    assign memory1a[19  ] = 3'd0;
    assign memory1a[20  ] = 3'd0;
    assign memory1a[21  ] = 3'd0;
    assign memory1a[22  ] = 3'd1;
    assign memory1a[23  ] = 3'd1;
    assign memory1a[24  ] = 3'd0;
    assign memory1a[25  ] = 3'd0;
    assign memory1a[26  ] = 3'd0;
    assign memory1a[27  ] = 3'd0;
    assign memory1a[28  ] = 3'd0;
    assign memory1a[29  ] = 3'd0;
    assign memory1a[30  ] = 3'd0;
    assign memory1a[31  ] = 3'd0;
    assign memory1a[32  ] = 3'd0;
    assign memory1a[33  ] = 3'd2;
    assign memory1a[34  ] = 3'd2;
    assign memory1a[35  ] = 3'd2;
    assign memory1a[36  ] = 3'd2;
    assign memory1a[37  ] = 3'd2;
    assign memory1a[38  ] = 3'd2;
    assign memory1a[39  ] = 3'd2;
    assign memory1a[40  ] = 3'd2;
    assign memory1a[41  ] = 3'd2;
    assign memory1a[42  ] = 3'd2;
    assign memory1a[43  ] = 3'd2;
    assign memory1a[44  ] = 3'd2;
    assign memory1a[45  ] = 3'd3;
    assign memory1a[46  ] = 3'd3;
    assign memory1a[47  ] = 3'd3;
    assign memory1a[48  ] = 3'd3;
    assign memory1a[49  ] = 3'd3;
    assign memory1a[50  ] = 3'd3;
    assign memory1a[51  ] = 3'd3;
    assign memory1a[52  ] = 3'd3;
    assign memory1a[53  ] = 3'd2;
    assign memory1a[54  ] = 3'd2;
    assign memory1a[55  ] = 3'd2;
    assign memory1a[56  ] = 3'd2;
    assign memory1a[57  ] = 3'd2;
    assign memory1a[58  ] = 3'd2;
    assign memory1a[59  ] = 3'd2;
    assign memory1a[60  ] = 3'd3;
    assign memory1a[61  ] = 3'd3;
    assign memory1a[62  ] = 3'd3;
    assign memory1a[63  ] = 3'd0;
    assign memory1a[64  ] = 3'd0;
    assign memory1a[65  ] = 3'd3;
    assign memory1a[66  ] = 3'd3;
    assign memory1a[67  ] = 3'd3;
    assign memory1a[68  ] = 3'd3;
    assign memory1a[69  ] = 3'd3;
    assign memory1a[70  ] = 3'd3;
    assign memory1a[71  ] = 3'd3;
    assign memory1a[72  ] = 3'd3;
    assign memory1a[73  ] = 3'd3;
    assign memory1a[74  ] = 3'd3;
    assign memory1a[75  ] = 3'd3;
    assign memory1a[76  ] = 3'd3;
    assign memory1a[77  ] = 3'd3;
    assign memory1a[78  ] = 3'd3;
    assign memory1a[79  ] = 3'd4;
    assign memory1a[80  ] = 3'd4;
    assign memory1a[81  ] = 3'd4;
    assign memory1a[82  ] = 3'd4;
    assign memory1a[83  ] = 3'd4;
    assign memory1a[84  ] = 3'd3;
    assign memory1a[85  ] = 3'd3;
    assign memory1a[86  ] = 3'd3;
    assign memory1a[87  ] = 3'd3;
    assign memory1a[88  ] = 3'd3;
    assign memory1a[89  ] = 3'd3;
    assign memory1a[90  ] = 3'd3;
    assign memory1a[91  ] = 3'd3;
    assign memory1a[92  ] = 3'd3;
    assign memory1a[93  ] = 3'd4;
    assign memory1a[94  ] = 3'd5;
    assign memory1a[95  ] = 3'd0;
    assign memory1a[96  ] = 3'd0;
    assign memory1a[97  ] = 3'd3;
    assign memory1a[98  ] = 3'd3;
    assign memory1a[99  ] = 3'd3;
    assign memory1a[100 ] = 3'd3;
    assign memory1a[101 ] = 3'd3;
    assign memory1a[102 ] = 3'd3;
    assign memory1a[103 ] = 3'd3;
    assign memory1a[104 ] = 3'd3;
    assign memory1a[105 ] = 3'd3;
    assign memory1a[106 ] = 3'd3;
    assign memory1a[107 ] = 3'd4;
    assign memory1a[108 ] = 3'd4;
    assign memory1a[109 ] = 3'd4;
    assign memory1a[110 ] = 3'd4;
    assign memory1a[111 ] = 3'd4;
    assign memory1a[112 ] = 3'd4;
    assign memory1a[113 ] = 3'd4;
    assign memory1a[114 ] = 3'd4;
    assign memory1a[115 ] = 3'd4;
    assign memory1a[116 ] = 3'd4;
    assign memory1a[117 ] = 3'd4;
    assign memory1a[118 ] = 3'd4;
    assign memory1a[119 ] = 3'd4;
    assign memory1a[120 ] = 3'd4;
    assign memory1a[121 ] = 3'd4;
    assign memory1a[122 ] = 3'd5;
    assign memory1a[123 ] = 3'd5;
    assign memory1a[124 ] = 3'd4;
    assign memory1a[125 ] = 3'd4;
    assign memory1a[126 ] = 3'd5;
    assign memory1a[127 ] = 3'd0;
    assign memory1a[128 ] = 3'd0;
    assign memory1a[129 ] = 3'd3;
    assign memory1a[130 ] = 3'd3;
    assign memory1a[131 ] = 3'd4;
    assign memory1a[132 ] = 3'd4;
    assign memory1a[133 ] = 3'd4;
    assign memory1a[134 ] = 3'd4;
    assign memory1a[135 ] = 3'd4;
    assign memory1a[136 ] = 3'd4;
    assign memory1a[137 ] = 3'd4;
    assign memory1a[138 ] = 3'd4;
    assign memory1a[139 ] = 3'd4;
    assign memory1a[140 ] = 3'd4;
    assign memory1a[141 ] = 3'd4;
    assign memory1a[142 ] = 3'd5;
    assign memory1a[143 ] = 3'd5;
    assign memory1a[144 ] = 3'd4;
    assign memory1a[145 ] = 3'd4;
    assign memory1a[146 ] = 3'd4;
    assign memory1a[147 ] = 3'd4;
    assign memory1a[148 ] = 3'd4;
    assign memory1a[149 ] = 3'd4;
    assign memory1a[150 ] = 3'd4;
    assign memory1a[151 ] = 3'd4;
    assign memory1a[152 ] = 3'd5;
    assign memory1a[153 ] = 3'd5;
    assign memory1a[154 ] = 3'd5;
    assign memory1a[155 ] = 3'd5;
    assign memory1a[156 ] = 3'd4;
    assign memory1a[157 ] = 3'd4;
    assign memory1a[158 ] = 3'd5;
    assign memory1a[159 ] = 3'd0;
    assign memory1a[160 ] = 3'd0;
    assign memory1a[161 ] = 3'd3;
    assign memory1a[162 ] = 3'd3;
    assign memory1a[163 ] = 3'd4;
    assign memory1a[164 ] = 3'd4;
    assign memory1a[165 ] = 3'd4;
    assign memory1a[166 ] = 3'd4;
    assign memory1a[167 ] = 3'd5;
    assign memory1a[168 ] = 3'd4;
    assign memory1a[169 ] = 3'd4;
    assign memory1a[170 ] = 3'd4;
    assign memory1a[171 ] = 3'd4;
    assign memory1a[172 ] = 3'd4;
    assign memory1a[173 ] = 3'd4;
    assign memory1a[174 ] = 3'd5;
    assign memory1a[175 ] = 3'd5;
    assign memory1a[176 ] = 3'd5;
    assign memory1a[177 ] = 3'd5;
    assign memory1a[178 ] = 3'd4;
    assign memory1a[179 ] = 3'd4;
    assign memory1a[180 ] = 3'd4;
    assign memory1a[181 ] = 3'd4;
    assign memory1a[182 ] = 3'd4;
    assign memory1a[183 ] = 3'd4;
    assign memory1a[184 ] = 3'd4;
    assign memory1a[185 ] = 3'd5;
    assign memory1a[186 ] = 3'd5;
    assign memory1a[187 ] = 3'd5;
    assign memory1a[188 ] = 3'd4;
    assign memory1a[189 ] = 3'd4;
    assign memory1a[190 ] = 3'd5;
    assign memory1a[191 ] = 3'd0;
    assign memory1a[192 ] = 3'd1;
    assign memory1a[193 ] = 3'd2;
    assign memory1a[194 ] = 3'd3;
    assign memory1a[195 ] = 3'd4;
    assign memory1a[196 ] = 3'd4;
    assign memory1a[197 ] = 3'd4;
    assign memory1a[198 ] = 3'd5;
    assign memory1a[199 ] = 3'd5;
    assign memory1a[200 ] = 3'd5;
    assign memory1a[201 ] = 3'd5;
    assign memory1a[202 ] = 3'd5;
    assign memory1a[203 ] = 3'd4;
    assign memory1a[204 ] = 3'd4;
    assign memory1a[205 ] = 3'd4;
    assign memory1a[206 ] = 3'd4;
    assign memory1a[207 ] = 3'd4;
    assign memory1a[208 ] = 3'd4;
    assign memory1a[209 ] = 3'd4;
    assign memory1a[210 ] = 3'd4;
    assign memory1a[211 ] = 3'd4;
    assign memory1a[212 ] = 3'd4;
    assign memory1a[213 ] = 3'd4;
    assign memory1a[214 ] = 3'd4;
    assign memory1a[215 ] = 3'd4;
    assign memory1a[216 ] = 3'd4;
    assign memory1a[217 ] = 3'd4;
    assign memory1a[218 ] = 3'd5;
    assign memory1a[219 ] = 3'd5;
    assign memory1a[220 ] = 3'd4;
    assign memory1a[221 ] = 3'd4;
    assign memory1a[222 ] = 3'd5;
    assign memory1a[223 ] = 3'd1;
    assign memory1a[224 ] = 3'd1;
    assign memory1a[225 ] = 3'd2;
    assign memory1a[226 ] = 3'd3;
    assign memory1a[227 ] = 3'd4;
    assign memory1a[228 ] = 3'd4;
    assign memory1a[229 ] = 3'd4;
    assign memory1a[230 ] = 3'd5;
    assign memory1a[231 ] = 3'd5;
    assign memory1a[232 ] = 3'd4;
    assign memory1a[233 ] = 3'd5;
    assign memory1a[234 ] = 3'd4;
    assign memory1a[235 ] = 3'd4;
    assign memory1a[236 ] = 3'd4;
    assign memory1a[237 ] = 3'd4;
    assign memory1a[238 ] = 3'd4;
    assign memory1a[239 ] = 3'd4;
    assign memory1a[240 ] = 3'd4;
    assign memory1a[241 ] = 3'd4;
    assign memory1a[242 ] = 3'd4;
    assign memory1a[243 ] = 3'd4;
    assign memory1a[244 ] = 3'd4;
    assign memory1a[245 ] = 3'd4;
    assign memory1a[246 ] = 3'd4;
    assign memory1a[247 ] = 3'd4;
    assign memory1a[248 ] = 3'd4;
    assign memory1a[249 ] = 3'd4;
    assign memory1a[250 ] = 3'd4;
    assign memory1a[251 ] = 3'd4;
    assign memory1a[252 ] = 3'd4;
    assign memory1a[253 ] = 3'd4;
    assign memory1a[254 ] = 3'd5;
    assign memory1a[255 ] = 3'd1;
    assign memory1a[256 ] = 3'd0;
    assign memory1a[257 ] = 3'd2;
    assign memory1a[258 ] = 3'd3;
    assign memory1a[259 ] = 3'd4;
    assign memory1a[260 ] = 3'd4;
    assign memory1a[261 ] = 3'd4;
    assign memory1a[262 ] = 3'd4;
    assign memory1a[263 ] = 3'd4;
    assign memory1a[264 ] = 3'd4;
    assign memory1a[265 ] = 3'd4;
    assign memory1a[266 ] = 3'd4;
    assign memory1a[267 ] = 3'd4;
    assign memory1a[268 ] = 3'd4;
    assign memory1a[269 ] = 3'd4;
    assign memory1a[270 ] = 3'd4;
    assign memory1a[271 ] = 3'd4;
    assign memory1a[272 ] = 3'd4;
    assign memory1a[273 ] = 3'd4;
    assign memory1a[274 ] = 3'd4;
    assign memory1a[275 ] = 3'd4;
    assign memory1a[276 ] = 3'd4;
    assign memory1a[277 ] = 3'd4;
    assign memory1a[278 ] = 3'd4;
    assign memory1a[279 ] = 3'd4;
    assign memory1a[280 ] = 3'd4;
    assign memory1a[281 ] = 3'd4;
    assign memory1a[282 ] = 3'd4;
    assign memory1a[283 ] = 3'd4;
    assign memory1a[284 ] = 3'd4;
    assign memory1a[285 ] = 3'd4;
    assign memory1a[286 ] = 3'd5;
    assign memory1a[287 ] = 3'd0;
    assign memory1a[288 ] = 3'd0;
    assign memory1a[289 ] = 3'd2;
    assign memory1a[290 ] = 3'd3;
    assign memory1a[291 ] = 3'd6;
    assign memory1a[292 ] = 3'd6;
    assign memory1a[293 ] = 3'd6;
    assign memory1a[294 ] = 3'd6;
    assign memory1a[295 ] = 3'd4;
    assign memory1a[296 ] = 3'd4;
    assign memory1a[297 ] = 3'd4;
    assign memory1a[298 ] = 3'd4;
    assign memory1a[299 ] = 3'd4;
    assign memory1a[300 ] = 3'd4;
    assign memory1a[301 ] = 3'd6;
    assign memory1a[302 ] = 3'd6;
    assign memory1a[303 ] = 3'd6;
    assign memory1a[304 ] = 3'd6;
    assign memory1a[305 ] = 3'd6;
    assign memory1a[306 ] = 3'd6;
    assign memory1a[307 ] = 3'd6;
    assign memory1a[308 ] = 3'd6;
    assign memory1a[309 ] = 3'd6;
    assign memory1a[310 ] = 3'd6;
    assign memory1a[311 ] = 3'd6;
    assign memory1a[312 ] = 3'd6;
    assign memory1a[313 ] = 3'd6;
    assign memory1a[314 ] = 3'd6;
    assign memory1a[315 ] = 3'd6;
    assign memory1a[316 ] = 3'd6;
    assign memory1a[317 ] = 3'd6;
    assign memory1a[318 ] = 3'd5;
    assign memory1a[319 ] = 3'd0;
    assign memory1a[320 ] = 3'd0;
    assign memory1a[321 ] = 3'd2;
    assign memory1a[322 ] = 3'd3;
    assign memory1a[323 ] = 3'd6;
    assign memory1a[324 ] = 3'd6;
    assign memory1a[325 ] = 3'd6;
    assign memory1a[326 ] = 3'd6;
    assign memory1a[327 ] = 3'd6;
    assign memory1a[328 ] = 3'd6;
    assign memory1a[329 ] = 3'd6;
    assign memory1a[330 ] = 3'd6;
    assign memory1a[331 ] = 3'd6;
    assign memory1a[332 ] = 3'd6;
    assign memory1a[333 ] = 3'd6;
    assign memory1a[334 ] = 3'd6;
    assign memory1a[335 ] = 3'd6;
    assign memory1a[336 ] = 3'd6;
    assign memory1a[337 ] = 3'd6;
    assign memory1a[338 ] = 3'd6;
    assign memory1a[339 ] = 3'd6;
    assign memory1a[340 ] = 3'd6;
    assign memory1a[341 ] = 3'd6;
    assign memory1a[342 ] = 3'd6;
    assign memory1a[343 ] = 3'd6;
    assign memory1a[344 ] = 3'd6;
    assign memory1a[345 ] = 3'd6;
    assign memory1a[346 ] = 3'd6;
    assign memory1a[347 ] = 3'd6;
    assign memory1a[348 ] = 3'd6;
    assign memory1a[349 ] = 3'd6;
    assign memory1a[350 ] = 3'd5;
    assign memory1a[351 ] = 3'd0;
    assign memory1a[352 ] = 3'd0;
    assign memory1a[353 ] = 3'd2;
    assign memory1a[354 ] = 3'd3;
    assign memory1a[355 ] = 3'd6;
    assign memory1a[356 ] = 3'd5;
    assign memory1a[357 ] = 3'd5;
    assign memory1a[358 ] = 3'd6;
    assign memory1a[359 ] = 3'd6;
    assign memory1a[360 ] = 3'd6;
    assign memory1a[361 ] = 3'd6;
    assign memory1a[362 ] = 3'd6;
    assign memory1a[363 ] = 3'd6;
    assign memory1a[364 ] = 3'd6;
    assign memory1a[365 ] = 3'd6;
    assign memory1a[366 ] = 3'd6;
    assign memory1a[367 ] = 3'd6;
    assign memory1a[368 ] = 3'd6;
    assign memory1a[369 ] = 3'd6;
    assign memory1a[370 ] = 3'd6;
    assign memory1a[371 ] = 3'd6;
    assign memory1a[372 ] = 3'd6;
    assign memory1a[373 ] = 3'd6;
    assign memory1a[374 ] = 3'd6;
    assign memory1a[375 ] = 3'd6;
    assign memory1a[376 ] = 3'd5;
    assign memory1a[377 ] = 3'd5;
    assign memory1a[378 ] = 3'd5;
    assign memory1a[379 ] = 3'd6;
    assign memory1a[380 ] = 3'd6;
    assign memory1a[381 ] = 3'd6;
    assign memory1a[382 ] = 3'd5;
    assign memory1a[383 ] = 3'd0;
    assign memory1a[384 ] = 3'd0;
    assign memory1a[385 ] = 3'd3;
    assign memory1a[386 ] = 3'd3;
    assign memory1a[387 ] = 3'd6;
    assign memory1a[388 ] = 3'd5;
    assign memory1a[389 ] = 3'd5;
    assign memory1a[390 ] = 3'd5;
    assign memory1a[391 ] = 3'd5;
    assign memory1a[392 ] = 3'd5;
    assign memory1a[393 ] = 3'd6;
    assign memory1a[394 ] = 3'd6;
    assign memory1a[395 ] = 3'd6;
    assign memory1a[396 ] = 3'd6;
    assign memory1a[397 ] = 3'd5;
    assign memory1a[398 ] = 3'd5;
    assign memory1a[399 ] = 3'd6;
    assign memory1a[400 ] = 3'd6;
    assign memory1a[401 ] = 3'd5;
    assign memory1a[402 ] = 3'd5;
    assign memory1a[403 ] = 3'd5;
    assign memory1a[404 ] = 3'd6;
    assign memory1a[405 ] = 3'd6;
    assign memory1a[406 ] = 3'd6;
    assign memory1a[407 ] = 3'd5;
    assign memory1a[408 ] = 3'd5;
    assign memory1a[409 ] = 3'd5;
    assign memory1a[410 ] = 3'd5;
    assign memory1a[411 ] = 3'd6;
    assign memory1a[412 ] = 3'd5;
    assign memory1a[413 ] = 3'd5;
    assign memory1a[414 ] = 3'd5;
    assign memory1a[415 ] = 3'd0;
    assign memory1a[416 ] = 3'd1;
    assign memory1a[417 ] = 3'd3;
    assign memory1a[418 ] = 3'd3;
    assign memory1a[419 ] = 3'd6;
    assign memory1a[420 ] = 3'd5;
    assign memory1a[421 ] = 3'd5;
    assign memory1a[422 ] = 3'd5;
    assign memory1a[423 ] = 3'd5;
    assign memory1a[424 ] = 3'd5;
    assign memory1a[425 ] = 3'd5;
    assign memory1a[426 ] = 3'd5;
    assign memory1a[427 ] = 3'd5;
    assign memory1a[428 ] = 3'd5;
    assign memory1a[429 ] = 3'd5;
    assign memory1a[430 ] = 3'd5;
    assign memory1a[431 ] = 3'd5;
    assign memory1a[432 ] = 3'd5;
    assign memory1a[433 ] = 3'd5;
    assign memory1a[434 ] = 3'd5;
    assign memory1a[435 ] = 3'd5;
    assign memory1a[436 ] = 3'd5;
    assign memory1a[437 ] = 3'd5;
    assign memory1a[438 ] = 3'd6;
    assign memory1a[439 ] = 3'd5;
    assign memory1a[440 ] = 3'd5;
    assign memory1a[441 ] = 3'd5;
    assign memory1a[442 ] = 3'd5;
    assign memory1a[443 ] = 3'd5;
    assign memory1a[444 ] = 3'd5;
    assign memory1a[445 ] = 3'd5;
    assign memory1a[446 ] = 3'd5;
    assign memory1a[447 ] = 3'd1;
    assign memory1a[448 ] = 3'd0;
    assign memory1a[449 ] = 3'd3;
    assign memory1a[450 ] = 3'd3;
    assign memory1a[451 ] = 3'd5;
    assign memory1a[452 ] = 3'd5;
    assign memory1a[453 ] = 3'd5;
    assign memory1a[454 ] = 3'd5;
    assign memory1a[455 ] = 3'd5;
    assign memory1a[456 ] = 3'd5;
    assign memory1a[457 ] = 3'd5;
    assign memory1a[458 ] = 3'd5;
    assign memory1a[459 ] = 3'd5;
    assign memory1a[460 ] = 3'd5;
    assign memory1a[461 ] = 3'd5;
    assign memory1a[462 ] = 3'd5;
    assign memory1a[463 ] = 3'd5;
    assign memory1a[464 ] = 3'd5;
    assign memory1a[465 ] = 3'd5;
    assign memory1a[466 ] = 3'd5;
    assign memory1a[467 ] = 3'd5;
    assign memory1a[468 ] = 3'd5;
    assign memory1a[469 ] = 3'd5;
    assign memory1a[470 ] = 3'd5;
    assign memory1a[471 ] = 3'd5;
    assign memory1a[472 ] = 3'd5;
    assign memory1a[473 ] = 3'd5;
    assign memory1a[474 ] = 3'd5;
    assign memory1a[475 ] = 3'd5;
    assign memory1a[476 ] = 3'd0;
    assign memory1a[477 ] = 3'd0;
    assign memory1a[478 ] = 3'd0;
    assign memory1a[479 ] = 3'd0;
    assign memory1a[480 ] = 3'd0;
    assign memory1a[481 ] = 3'd0;
    assign memory1a[482 ] = 3'd0;
    assign memory1a[483 ] = 3'd0;
    assign memory1a[484 ] = 3'd0;
    assign memory1a[485 ] = 3'd0;
    assign memory1a[486 ] = 3'd0;
    assign memory1a[487 ] = 3'd0;
    assign memory1a[488 ] = 3'd0;
    assign memory1a[489 ] = 3'd0;
    assign memory1a[490 ] = 3'd1;
    assign memory1a[491 ] = 3'd0;
    assign memory1a[492 ] = 3'd0;
    assign memory1a[493 ] = 3'd0;
    assign memory1a[494 ] = 3'd0;
    assign memory1a[495 ] = 3'd0;
    assign memory1a[496 ] = 3'd0;
    assign memory1a[497 ] = 3'd0;
    assign memory1a[498 ] = 3'd0;
    assign memory1a[499 ] = 3'd0;
    assign memory1a[500 ] = 3'd0;
    assign memory1a[501 ] = 3'd0;
    assign memory1a[502 ] = 3'd0;
    assign memory1a[503 ] = 3'd0;
    assign memory1a[504 ] = 3'd0;
    assign memory1a[505 ] = 3'd1;
    assign memory1a[506 ] = 3'd1;
    assign memory1a[507 ] = 3'd0;
    assign memory1a[508 ] = 3'd0;
    assign memory1a[509 ] = 3'd0;
    assign memory1a[510 ] = 3'd0;
    assign memory1a[511 ] = 3'd0;
    assign memory1a[512 ] = 3'd0;
    assign memory1a[513 ] = 3'd0;
    assign memory1a[514 ] = 3'd0;
    assign memory1a[515 ] = 3'd0;
    assign memory1a[516 ] = 3'd0;
    assign memory1a[517 ] = 3'd0;
    assign memory1a[518 ] = 3'd0;
    assign memory1a[519 ] = 3'd0;
    assign memory1a[520 ] = 3'd0;
    assign memory1a[521 ] = 3'd0;
    assign memory1a[522 ] = 3'd1;
    assign memory1a[523 ] = 3'd0;
    assign memory1a[524 ] = 3'd0;
    assign memory1a[525 ] = 3'd0;
    assign memory1a[526 ] = 3'd0;
    assign memory1a[527 ] = 3'd0;
    assign memory1a[528 ] = 3'd0;
    assign memory1a[529 ] = 3'd0;
    assign memory1a[530 ] = 3'd0;
    assign memory1a[531 ] = 3'd0;
    assign memory1a[532 ] = 3'd0;
    assign memory1a[533 ] = 3'd0;
    assign memory1a[534 ] = 3'd0;
    assign memory1a[535 ] = 3'd0;
    assign memory1a[536 ] = 3'd0;
    assign memory1a[537 ] = 3'd1;
    assign memory1a[538 ] = 3'd1;
    assign memory1a[539 ] = 3'd0;
    assign memory1a[540 ] = 3'd0;
    assign memory1a[541 ] = 3'd0;
    assign memory1a[542 ] = 3'd0;
    assign memory1a[543 ] = 3'd0;
    assign memory1a[544 ] = 3'd3;
    assign memory1a[545 ] = 3'd3;
    assign memory1a[546 ] = 3'd3;
    assign memory1a[547 ] = 3'd3;
    assign memory1a[548 ] = 3'd3;
    assign memory1a[549 ] = 3'd3;
    assign memory1a[550 ] = 3'd3;
    assign memory1a[551 ] = 3'd3;
    assign memory1a[552 ] = 3'd3;
    assign memory1a[553 ] = 3'd3;
    assign memory1a[554 ] = 3'd3;
    assign memory1a[555 ] = 3'd3;
    assign memory1a[556 ] = 3'd3;
    assign memory1a[557 ] = 3'd3;
    assign memory1a[558 ] = 3'd2;
    assign memory1a[559 ] = 3'd0;
    assign memory1a[560 ] = 3'd0;
    assign memory1a[561 ] = 3'd2;
    assign memory1a[562 ] = 3'd2;
    assign memory1a[563 ] = 3'd3;
    assign memory1a[564 ] = 3'd3;
    assign memory1a[565 ] = 3'd3;
    assign memory1a[566 ] = 3'd3;
    assign memory1a[567 ] = 3'd3;
    assign memory1a[568 ] = 3'd3;
    assign memory1a[569 ] = 3'd3;
    assign memory1a[570 ] = 3'd3;
    assign memory1a[571 ] = 3'd3;
    assign memory1a[572 ] = 3'd3;
    assign memory1a[573 ] = 3'd3;
    assign memory1a[574 ] = 3'd3;
    assign memory1a[575 ] = 3'd3;
    assign memory1a[576 ] = 3'd3;
    assign memory1a[577 ] = 3'd4;
    assign memory1a[578 ] = 3'd4;
    assign memory1a[579 ] = 3'd4;
    assign memory1a[580 ] = 3'd4;
    assign memory1a[581 ] = 3'd4;
    assign memory1a[582 ] = 3'd4;
    assign memory1a[583 ] = 3'd4;
    assign memory1a[584 ] = 3'd4;
    assign memory1a[585 ] = 3'd4;
    assign memory1a[586 ] = 3'd4;
    assign memory1a[587 ] = 3'd4;
    assign memory1a[588 ] = 3'd4;
    assign memory1a[589 ] = 3'd4;
    assign memory1a[590 ] = 3'd5;
    assign memory1a[591 ] = 3'd0;
    assign memory1a[592 ] = 3'd0;
    assign memory1a[593 ] = 3'd3;
    assign memory1a[594 ] = 3'd3;
    assign memory1a[595 ] = 3'd3;
    assign memory1a[596 ] = 3'd3;
    assign memory1a[597 ] = 3'd3;
    assign memory1a[598 ] = 3'd3;
    assign memory1a[599 ] = 3'd3;
    assign memory1a[600 ] = 3'd3;
    assign memory1a[601 ] = 3'd3;
    assign memory1a[602 ] = 3'd3;
    assign memory1a[603 ] = 3'd3;
    assign memory1a[604 ] = 3'd3;
    assign memory1a[605 ] = 3'd3;
    assign memory1a[606 ] = 3'd3;
    assign memory1a[607 ] = 3'd3;
    assign memory1a[608 ] = 3'd4;
    assign memory1a[609 ] = 3'd4;
    assign memory1a[610 ] = 3'd4;
    assign memory1a[611 ] = 3'd4;
    assign memory1a[612 ] = 3'd4;
    assign memory1a[613 ] = 3'd4;
    assign memory1a[614 ] = 3'd4;
    assign memory1a[615 ] = 3'd4;
    assign memory1a[616 ] = 3'd4;
    assign memory1a[617 ] = 3'd5;
    assign memory1a[618 ] = 3'd4;
    assign memory1a[619 ] = 3'd4;
    assign memory1a[620 ] = 3'd4;
    assign memory1a[621 ] = 3'd4;
    assign memory1a[622 ] = 3'd5;
    assign memory1a[623 ] = 3'd0;
    assign memory1a[624 ] = 3'd0;
    assign memory1a[625 ] = 3'd3;
    assign memory1a[626 ] = 3'd3;
    assign memory1a[627 ] = 3'd4;
    assign memory1a[628 ] = 3'd4;
    assign memory1a[629 ] = 3'd4;
    assign memory1a[630 ] = 3'd4;
    assign memory1a[631 ] = 3'd4;
    assign memory1a[632 ] = 3'd4;
    assign memory1a[633 ] = 3'd4;
    assign memory1a[634 ] = 3'd4;
    assign memory1a[635 ] = 3'd4;
    assign memory1a[636 ] = 3'd4;
    assign memory1a[637 ] = 3'd4;
    assign memory1a[638 ] = 3'd4;
    assign memory1a[639 ] = 3'd4;
    assign memory1a[640 ] = 3'd4;
    assign memory1a[641 ] = 3'd4;
    assign memory1a[642 ] = 3'd4;
    assign memory1a[643 ] = 3'd4;
    assign memory1a[644 ] = 3'd4;
    assign memory1a[645 ] = 3'd4;
    assign memory1a[646 ] = 3'd5;
    assign memory1a[647 ] = 3'd5;
    assign memory1a[648 ] = 3'd5;
    assign memory1a[649 ] = 3'd5;
    assign memory1a[650 ] = 3'd5;
    assign memory1a[651 ] = 3'd4;
    assign memory1a[652 ] = 3'd4;
    assign memory1a[653 ] = 3'd4;
    assign memory1a[654 ] = 3'd5;
    assign memory1a[655 ] = 3'd1;
    assign memory1a[656 ] = 3'd1;
    assign memory1a[657 ] = 3'd3;
    assign memory1a[658 ] = 3'd3;
    assign memory1a[659 ] = 3'd4;
    assign memory1a[660 ] = 3'd4;
    assign memory1a[661 ] = 3'd4;
    assign memory1a[662 ] = 3'd4;
    assign memory1a[663 ] = 3'd4;
    assign memory1a[664 ] = 3'd4;
    assign memory1a[665 ] = 3'd5;
    assign memory1a[666 ] = 3'd4;
    assign memory1a[667 ] = 3'd4;
    assign memory1a[668 ] = 3'd4;
    assign memory1a[669 ] = 3'd4;
    assign memory1a[670 ] = 3'd4;
    assign memory1a[671 ] = 3'd4;
    assign memory1a[672 ] = 3'd5;
    assign memory1a[673 ] = 3'd5;
    assign memory1a[674 ] = 3'd4;
    assign memory1a[675 ] = 3'd4;
    assign memory1a[676 ] = 3'd4;
    assign memory1a[677 ] = 3'd4;
    assign memory1a[678 ] = 3'd4;
    assign memory1a[679 ] = 3'd4;
    assign memory1a[680 ] = 3'd5;
    assign memory1a[681 ] = 3'd5;
    assign memory1a[682 ] = 3'd5;
    assign memory1a[683 ] = 3'd4;
    assign memory1a[684 ] = 3'd4;
    assign memory1a[685 ] = 3'd4;
    assign memory1a[686 ] = 3'd5;
    assign memory1a[687 ] = 3'd1;
    assign memory1a[688 ] = 3'd1;
    assign memory1a[689 ] = 3'd3;
    assign memory1a[690 ] = 3'd3;
    assign memory1a[691 ] = 3'd4;
    assign memory1a[692 ] = 3'd5;
    assign memory1a[693 ] = 3'd5;
    assign memory1a[694 ] = 3'd4;
    assign memory1a[695 ] = 3'd4;
    assign memory1a[696 ] = 3'd4;
    assign memory1a[697 ] = 3'd4;
    assign memory1a[698 ] = 3'd4;
    assign memory1a[699 ] = 3'd4;
    assign memory1a[700 ] = 3'd4;
    assign memory1a[701 ] = 3'd5;
    assign memory1a[702 ] = 3'd5;
    assign memory1a[703 ] = 3'd5;
    assign memory1a[704 ] = 3'd5;
    assign memory1a[705 ] = 3'd5;
    assign memory1a[706 ] = 3'd4;
    assign memory1a[707 ] = 3'd4;
    assign memory1a[708 ] = 3'd4;
    assign memory1a[709 ] = 3'd4;
    assign memory1a[710 ] = 3'd4;
    assign memory1a[711 ] = 3'd4;
    assign memory1a[712 ] = 3'd4;
    assign memory1a[713 ] = 3'd4;
    assign memory1a[714 ] = 3'd4;
    assign memory1a[715 ] = 3'd4;
    assign memory1a[716 ] = 3'd4;
    assign memory1a[717 ] = 3'd4;
    assign memory1a[718 ] = 3'd5;
    assign memory1a[719 ] = 3'd0;
    assign memory1a[720 ] = 3'd0;
    assign memory1a[721 ] = 3'd3;
    assign memory1a[722 ] = 3'd3;
    assign memory1a[723 ] = 3'd4;
    assign memory1a[724 ] = 3'd5;
    assign memory1a[725 ] = 3'd5;
    assign memory1a[726 ] = 3'd5;
    assign memory1a[727 ] = 3'd4;
    assign memory1a[728 ] = 3'd4;
    assign memory1a[729 ] = 3'd4;
    assign memory1a[730 ] = 3'd4;
    assign memory1a[731 ] = 3'd4;
    assign memory1a[732 ] = 3'd4;
    assign memory1a[733 ] = 3'd4;
    assign memory1a[734 ] = 3'd5;
    assign memory1a[735 ] = 3'd5;
    assign memory1a[736 ] = 3'd4;
    assign memory1a[737 ] = 3'd4;
    assign memory1a[738 ] = 3'd4;
    assign memory1a[739 ] = 3'd4;
    assign memory1a[740 ] = 3'd4;
    assign memory1a[741 ] = 3'd4;
    assign memory1a[742 ] = 3'd4;
    assign memory1a[743 ] = 3'd4;
    assign memory1a[744 ] = 3'd4;
    assign memory1a[745 ] = 3'd4;
    assign memory1a[746 ] = 3'd4;
    assign memory1a[747 ] = 3'd4;
    assign memory1a[748 ] = 3'd4;
    assign memory1a[749 ] = 3'd4;
    assign memory1a[750 ] = 3'd5;
    assign memory1a[751 ] = 3'd0;
    assign memory1a[752 ] = 3'd0;
    assign memory1a[753 ] = 3'd3;
    assign memory1a[754 ] = 3'd3;
    assign memory1a[755 ] = 3'd4;
    assign memory1a[756 ] = 3'd4;
    assign memory1a[757 ] = 3'd5;
    assign memory1a[758 ] = 3'd4;
    assign memory1a[759 ] = 3'd4;
    assign memory1a[760 ] = 3'd4;
    assign memory1a[761 ] = 3'd4;
    assign memory1a[762 ] = 3'd4;
    assign memory1a[763 ] = 3'd4;
    assign memory1a[764 ] = 3'd4;
    assign memory1a[765 ] = 3'd4;
    assign memory1a[766 ] = 3'd4;
    assign memory1a[767 ] = 3'd4;
    assign memory1a[768 ] = 3'd4;
    assign memory1a[769 ] = 3'd4;
    assign memory1a[770 ] = 3'd6;
    assign memory1a[771 ] = 3'd6;
    assign memory1a[772 ] = 3'd6;
    assign memory1a[773 ] = 3'd6;
    assign memory1a[774 ] = 3'd6;
    assign memory1a[775 ] = 3'd6;
    assign memory1a[776 ] = 3'd6;
    assign memory1a[777 ] = 3'd6;
    assign memory1a[778 ] = 3'd4;
    assign memory1a[779 ] = 3'd4;
    assign memory1a[780 ] = 3'd4;
    assign memory1a[781 ] = 3'd4;
    assign memory1a[782 ] = 3'd5;
    assign memory1a[783 ] = 3'd0;
    assign memory1a[784 ] = 3'd0;
    assign memory1a[785 ] = 3'd3;
    assign memory1a[786 ] = 3'd3;
    assign memory1a[787 ] = 3'd4;
    assign memory1a[788 ] = 3'd4;
    assign memory1a[789 ] = 3'd4;
    assign memory1a[790 ] = 3'd4;
    assign memory1a[791 ] = 3'd4;
    assign memory1a[792 ] = 3'd4;
    assign memory1a[793 ] = 3'd4;
    assign memory1a[794 ] = 3'd4;
    assign memory1a[795 ] = 3'd4;
    assign memory1a[796 ] = 3'd4;
    assign memory1a[797 ] = 3'd4;
    assign memory1a[798 ] = 3'd4;
    assign memory1a[799 ] = 3'd4;
    assign memory1a[800 ] = 3'd6;
    assign memory1a[801 ] = 3'd6;
    assign memory1a[802 ] = 3'd6;
    assign memory1a[803 ] = 3'd6;
    assign memory1a[804 ] = 3'd6;
    assign memory1a[805 ] = 3'd6;
    assign memory1a[806 ] = 3'd6;
    assign memory1a[807 ] = 3'd6;
    assign memory1a[808 ] = 3'd6;
    assign memory1a[809 ] = 3'd6;
    assign memory1a[810 ] = 3'd6;
    assign memory1a[811 ] = 3'd6;
    assign memory1a[812 ] = 3'd6;
    assign memory1a[813 ] = 3'd6;
    assign memory1a[814 ] = 3'd5;
    assign memory1a[815 ] = 3'd0;
    assign memory1a[816 ] = 3'd0;
    assign memory1a[817 ] = 3'd3;
    assign memory1a[818 ] = 3'd3;
    assign memory1a[819 ] = 3'd4;
    assign memory1a[820 ] = 3'd6;
    assign memory1a[821 ] = 3'd6;
    assign memory1a[822 ] = 3'd6;
    assign memory1a[823 ] = 3'd6;
    assign memory1a[824 ] = 3'd6;
    assign memory1a[825 ] = 3'd6;
    assign memory1a[826 ] = 3'd6;
    assign memory1a[827 ] = 3'd4;
    assign memory1a[828 ] = 3'd4;
    assign memory1a[829 ] = 3'd4;
    assign memory1a[830 ] = 3'd4;
    assign memory1a[831 ] = 3'd6;
    assign memory1a[832 ] = 3'd6;
    assign memory1a[833 ] = 3'd6;
    assign memory1a[834 ] = 3'd6;
    assign memory1a[835 ] = 3'd5;
    assign memory1a[836 ] = 3'd5;
    assign memory1a[837 ] = 3'd6;
    assign memory1a[838 ] = 3'd6;
    assign memory1a[839 ] = 3'd6;
    assign memory1a[840 ] = 3'd6;
    assign memory1a[841 ] = 3'd6;
    assign memory1a[842 ] = 3'd6;
    assign memory1a[843 ] = 3'd6;
    assign memory1a[844 ] = 3'd6;
    assign memory1a[845 ] = 3'd6;
    assign memory1a[846 ] = 3'd5;
    assign memory1a[847 ] = 3'd0;
    assign memory1a[848 ] = 3'd0;
    assign memory1a[849 ] = 3'd3;
    assign memory1a[850 ] = 3'd3;
    assign memory1a[851 ] = 3'd6;
    assign memory1a[852 ] = 3'd6;
    assign memory1a[853 ] = 3'd6;
    assign memory1a[854 ] = 3'd6;
    assign memory1a[855 ] = 3'd6;
    assign memory1a[856 ] = 3'd6;
    assign memory1a[857 ] = 3'd6;
    assign memory1a[858 ] = 3'd6;
    assign memory1a[859 ] = 3'd5;
    assign memory1a[860 ] = 3'd5;
    assign memory1a[861 ] = 3'd6;
    assign memory1a[862 ] = 3'd6;
    assign memory1a[863 ] = 3'd6;
    assign memory1a[864 ] = 3'd6;
    assign memory1a[865 ] = 3'd5;
    assign memory1a[866 ] = 3'd5;
    assign memory1a[867 ] = 3'd5;
    assign memory1a[868 ] = 3'd5;
    assign memory1a[869 ] = 3'd5;
    assign memory1a[870 ] = 3'd6;
    assign memory1a[871 ] = 3'd6;
    assign memory1a[872 ] = 3'd6;
    assign memory1a[873 ] = 3'd6;
    assign memory1a[874 ] = 3'd6;
    assign memory1a[875 ] = 3'd6;
    assign memory1a[876 ] = 3'd6;
    assign memory1a[877 ] = 3'd6;
    assign memory1a[878 ] = 3'd5;
    assign memory1a[879 ] = 3'd1;
    assign memory1a[880 ] = 3'd1;
    assign memory1a[881 ] = 3'd3;
    assign memory1a[882 ] = 3'd3;
    assign memory1a[883 ] = 3'd6;
    assign memory1a[884 ] = 3'd6;
    assign memory1a[885 ] = 3'd6;
    assign memory1a[886 ] = 3'd6;
    assign memory1a[887 ] = 3'd6;
    assign memory1a[888 ] = 3'd6;
    assign memory1a[889 ] = 3'd5;
    assign memory1a[890 ] = 3'd5;
    assign memory1a[891 ] = 3'd5;
    assign memory1a[892 ] = 3'd5;
    assign memory1a[893 ] = 3'd5;
    assign memory1a[894 ] = 3'd6;
    assign memory1a[895 ] = 3'd6;
    assign memory1a[896 ] = 3'd5;
    assign memory1a[897 ] = 3'd5;
    assign memory1a[898 ] = 3'd5;
    assign memory1a[899 ] = 3'd5;
    assign memory1a[900 ] = 3'd5;
    assign memory1a[901 ] = 3'd5;
    assign memory1a[902 ] = 3'd6;
    assign memory1a[903 ] = 3'd6;
    assign memory1a[904 ] = 3'd6;
    assign memory1a[905 ] = 3'd6;
    assign memory1a[906 ] = 3'd6;
    assign memory1a[907 ] = 3'd5;
    assign memory1a[908 ] = 3'd5;
    assign memory1a[909 ] = 3'd5;
    assign memory1a[910 ] = 3'd5;
    assign memory1a[911 ] = 3'd0;
    assign memory1a[912 ] = 3'd0;
    assign memory1a[913 ] = 3'd3;
    assign memory1a[914 ] = 3'd3;
    assign memory1a[915 ] = 3'd6;
    assign memory1a[916 ] = 3'd6;
    assign memory1a[917 ] = 3'd6;
    assign memory1a[918 ] = 3'd6;
    assign memory1a[919 ] = 3'd6;
    assign memory1a[920 ] = 3'd5;
    assign memory1a[921 ] = 3'd5;
    assign memory1a[922 ] = 3'd5;
    assign memory1a[923 ] = 3'd5;
    assign memory1a[924 ] = 3'd5;
    assign memory1a[925 ] = 3'd5;
    assign memory1a[926 ] = 3'd5;
    assign memory1a[927 ] = 3'd5;
    assign memory1a[928 ] = 3'd5;
    assign memory1a[929 ] = 3'd5;
    assign memory1a[930 ] = 3'd5;
    assign memory1a[931 ] = 3'd5;
    assign memory1a[932 ] = 3'd5;
    assign memory1a[933 ] = 3'd5;
    assign memory1a[934 ] = 3'd6;
    assign memory1a[935 ] = 3'd6;
    assign memory1a[936 ] = 3'd5;
    assign memory1a[937 ] = 3'd5;
    assign memory1a[938 ] = 3'd5;
    assign memory1a[939 ] = 3'd5;
    assign memory1a[940 ] = 3'd5;
    assign memory1a[941 ] = 3'd5;
    assign memory1a[942 ] = 3'd2;
    assign memory1a[943 ] = 3'd0;
    assign memory1a[944 ] = 3'd0;
    assign memory1a[945 ] = 3'd0;
    assign memory1a[946 ] = 3'd3;
    assign memory1a[947 ] = 3'd6;
    assign memory1a[948 ] = 3'd6;
    assign memory1a[949 ] = 3'd6;
    assign memory1a[950 ] = 3'd5;
    assign memory1a[951 ] = 3'd5;
    assign memory1a[952 ] = 3'd5;
    assign memory1a[953 ] = 3'd5;
    assign memory1a[954 ] = 3'd5;
    assign memory1a[955 ] = 3'd5;
    assign memory1a[956 ] = 3'd5;
    assign memory1a[957 ] = 3'd5;
    assign memory1a[958 ] = 3'd5;
    assign memory1a[959 ] = 3'd5;
    assign memory1a[960 ] = 3'd2;
    assign memory1a[961 ] = 3'd2;
    assign memory1a[962 ] = 3'd2;
    assign memory1a[963 ] = 3'd2;
    assign memory1a[964 ] = 3'd2;
    assign memory1a[965 ] = 3'd5;
    assign memory1a[966 ] = 3'd5;
    assign memory1a[967 ] = 3'd5;
    assign memory1a[968 ] = 3'd5;
    assign memory1a[969 ] = 3'd5;
    assign memory1a[970 ] = 3'd5;
    assign memory1a[971 ] = 3'd5;
    assign memory1a[972 ] = 3'd5;
    assign memory1a[973 ] = 3'd5;
    assign memory1a[974 ] = 3'd2;
    assign memory1a[975 ] = 3'd0;
    assign memory1a[976 ] = 3'd0;
    assign memory1a[977 ] = 3'd0;
    assign memory1a[978 ] = 3'd3;
    assign memory1a[979 ] = 3'd5;
    assign memory1a[980 ] = 3'd5;
    assign memory1a[981 ] = 3'd5;
    assign memory1a[982 ] = 3'd5;
    assign memory1a[983 ] = 3'd5;
    assign memory1a[984 ] = 3'd2;
    assign memory1a[985 ] = 3'd2;
    assign memory1a[986 ] = 3'd2;
    assign memory1a[987 ] = 3'd2;
    assign memory1a[988 ] = 3'd2;
    assign memory1a[989 ] = 3'd2;
    assign memory1a[990 ] = 3'd2;
    assign memory1a[991 ] = 3'd5;
    assign memory1a[992 ] = 3'd0;
    assign memory1a[993 ] = 3'd0;
    assign memory1a[994 ] = 3'd0;
    assign memory1a[995 ] = 3'd0;
    assign memory1a[996 ] = 3'd0;
    assign memory1a[997 ] = 3'd1;
    assign memory1a[998 ] = 3'd1;
    assign memory1a[999 ] = 3'd0;
    assign memory1a[1000] = 3'd0;
    assign memory1a[1001] = 3'd0;
    assign memory1a[1002] = 3'd0;
    assign memory1a[1003] = 3'd0;
    assign memory1a[1004] = 3'd0;
    assign memory1a[1005] = 3'd1;
    assign memory1a[1006] = 3'd0;
    assign memory1a[1007] = 3'd0;
    assign memory1a[1008] = 3'd0;
    assign memory1a[1009] = 3'd0;
    assign memory1a[1010] = 3'd0;
    assign memory1a[1011] = 3'd0;
    assign memory1a[1012] = 3'd0;
    assign memory1a[1013] = 3'd0;
    assign memory1a[1014] = 3'd1;
    assign memory1a[1015] = 3'd1;
    assign memory1a[1016] = 3'd0;
    assign memory1a[1017] = 3'd0;
    assign memory1a[1018] = 3'd0;
    assign memory1a[1019] = 3'd0;
    assign memory1a[1020] = 3'd0;
    assign memory1a[1021] = 3'd0;
    assign memory1a[1022] = 3'd0;
    assign memory1a[1023] = 3'd0;

    assign memory1b[0   ] = 3'd0;
    assign memory1b[1   ] = 3'd1;
    assign memory1b[2   ] = 3'd2;
    assign memory1b[3   ] = 3'd0;
    assign memory1b[4   ] = 3'd2;
    assign memory1b[5   ] = 3'd2;
    assign memory1b[6   ] = 3'd2;
    assign memory1b[7   ] = 3'd3;
    assign memory1b[8   ] = 3'd3;
    assign memory1b[9   ] = 3'd0;
    assign memory1b[10  ] = 3'd2;
    assign memory1b[11  ] = 3'd0;
    assign memory1b[12  ] = 3'd0;
    assign memory1b[13  ] = 3'd2;
    assign memory1b[14  ] = 3'd1;
    assign memory1b[15  ] = 3'd2;
    assign memory1b[16  ] = 3'd0;
    assign memory1b[17  ] = 3'd0;
    assign memory1b[18  ] = 3'd4;
    assign memory1b[19  ] = 3'd0;
    assign memory1b[20  ] = 3'd0;
    assign memory1b[21  ] = 3'd4;
    assign memory1b[22  ] = 3'd0;
    assign memory1b[23  ] = 3'd2;
    assign memory1b[24  ] = 3'd2;
    assign memory1b[25  ] = 3'd0;
    assign memory1b[26  ] = 3'd0;
    assign memory1b[27  ] = 3'd3;
    assign memory1b[28  ] = 3'd0;
    assign memory1b[29  ] = 3'd0;
    assign memory1b[30  ] = 3'd2;
    assign memory1b[31  ] = 3'd0;
    assign memory1b[32  ] = 3'd2;
    assign memory1b[33  ] = 3'd0;
    assign memory1b[34  ] = 3'd0;
    assign memory1b[35  ] = 3'd2;
    assign memory1b[36  ] = 3'd0;
    assign memory1b[37  ] = 3'd3;
    assign memory1b[38  ] = 3'd0;
    assign memory1b[39  ] = 3'd0;
    assign memory1b[40  ] = 3'd0;
    assign memory1b[41  ] = 3'd2;
    assign memory1b[42  ] = 3'd2;
    assign memory1b[43  ] = 3'd0;
    assign memory1b[44  ] = 3'd4;
    assign memory1b[45  ] = 3'd0;
    assign memory1b[46  ] = 3'd0;
    assign memory1b[47  ] = 3'd2;
    assign memory1b[48  ] = 3'd4;
    assign memory1b[49  ] = 3'd0;
    assign memory1b[50  ] = 3'd4;
    assign memory1b[51  ] = 3'd4;
    assign memory1b[52  ] = 3'd0;
    assign memory1b[53  ] = 3'd0;
    assign memory1b[54  ] = 3'd0;
    assign memory1b[55  ] = 3'd4;
    assign memory1b[56  ] = 3'd0;
    assign memory1b[57  ] = 3'd0;
    assign memory1b[58  ] = 3'd0;
    assign memory1b[59  ] = 3'd0;
    assign memory1b[60  ] = 3'd4;
    assign memory1b[61  ] = 3'd0;
    assign memory1b[62  ] = 3'd4;
    assign memory1b[63  ] = 3'd1;
    assign memory1b[64  ] = 3'd2;
    assign memory1b[65  ] = 3'd2;
    assign memory1b[66  ] = 3'd0;
    assign memory1b[67  ] = 3'd2;
    assign memory1b[68  ] = 3'd0;
    assign memory1b[69  ] = 3'd2;
    assign memory1b[70  ] = 3'd0;
    assign memory1b[71  ] = 3'd0;
    assign memory1b[72  ] = 3'd0;
    assign memory1b[73  ] = 3'd0;
    assign memory1b[74  ] = 3'd2;
    assign memory1b[75  ] = 3'd0;
    assign memory1b[76  ] = 3'd2;
    assign memory1b[77  ] = 3'd3;
    assign memory1b[78  ] = 3'd2;
    assign memory1b[79  ] = 3'd4;
    assign memory1b[80  ] = 3'd0;
    assign memory1b[81  ] = 3'd0;
    assign memory1b[82  ] = 3'd0;
    assign memory1b[83  ] = 3'd0;
    assign memory1b[84  ] = 3'd2;
    assign memory1b[85  ] = 3'd4;
    assign memory1b[86  ] = 3'd0;
    assign memory1b[87  ] = 3'd0;
    assign memory1b[88  ] = 3'd0;
    assign memory1b[89  ] = 3'd4;
    assign memory1b[90  ] = 3'd0;
    assign memory1b[91  ] = 3'd1;
    assign memory1b[92  ] = 3'd0;
    assign memory1b[93  ] = 3'd2;
    assign memory1b[94  ] = 3'd0;
    assign memory1b[95  ] = 3'd0;
    assign memory1b[96  ] = 3'd2;
    assign memory1b[97  ] = 3'd3;
    assign memory1b[98  ] = 3'd0;
    assign memory1b[99  ] = 3'd0;
    assign memory1b[100 ] = 3'd0;
    assign memory1b[101 ] = 3'd2;
    assign memory1b[102 ] = 3'd1;
    assign memory1b[103 ] = 3'd4;
    assign memory1b[104 ] = 3'd0;
    assign memory1b[105 ] = 3'd0;
    assign memory1b[106 ] = 3'd0;
    assign memory1b[107 ] = 3'd2;
    assign memory1b[108 ] = 3'd0;
    assign memory1b[109 ] = 3'd0;
    assign memory1b[110 ] = 3'd4;
    assign memory1b[111 ] = 3'd0;
    assign memory1b[112 ] = 3'd0;
    assign memory1b[113 ] = 3'd4;
    assign memory1b[114 ] = 3'd2;
    assign memory1b[115 ] = 3'd2;
    assign memory1b[116 ] = 3'd0;
    assign memory1b[117 ] = 3'd2;
    assign memory1b[118 ] = 3'd0;
    assign memory1b[119 ] = 3'd0;
    assign memory1b[120 ] = 3'd0;
    assign memory1b[121 ] = 3'd0;
    assign memory1b[122 ] = 3'd0;
    assign memory1b[123 ] = 3'd2;
    assign memory1b[124 ] = 3'd2;
    assign memory1b[125 ] = 3'd4;
    assign memory1b[126 ] = 3'd4;
    assign memory1b[127 ] = 3'd0;
    assign memory1b[128 ] = 3'd0;
    assign memory1b[129 ] = 3'd0;
    assign memory1b[130 ] = 3'd0;
    assign memory1b[131 ] = 3'd0;
    assign memory1b[132 ] = 3'd0;
    assign memory1b[133 ] = 3'd1;
    assign memory1b[134 ] = 3'd1;
    assign memory1b[135 ] = 3'd0;
    assign memory1b[136 ] = 3'd2;
    assign memory1b[137 ] = 3'd0;
    assign memory1b[138 ] = 3'd0;
    assign memory1b[139 ] = 3'd0;
    assign memory1b[140 ] = 3'd0;
    assign memory1b[141 ] = 3'd0;
    assign memory1b[142 ] = 3'd4;
    assign memory1b[143 ] = 3'd0;
    assign memory1b[144 ] = 3'd0;
    assign memory1b[145 ] = 3'd0;
    assign memory1b[146 ] = 3'd0;
    assign memory1b[147 ] = 3'd4;
    assign memory1b[148 ] = 3'd2;
    assign memory1b[149 ] = 3'd0;
    assign memory1b[150 ] = 3'd3;
    assign memory1b[151 ] = 3'd2;
    assign memory1b[152 ] = 3'd0;
    assign memory1b[153 ] = 3'd0;
    assign memory1b[154 ] = 3'd0;
    assign memory1b[155 ] = 3'd1;
    assign memory1b[156 ] = 3'd0;
    assign memory1b[157 ] = 3'd0;
    assign memory1b[158 ] = 3'd0;
    assign memory1b[159 ] = 3'd0;
    assign memory1b[160 ] = 3'd0;
    assign memory1b[161 ] = 3'd2;
    assign memory1b[162 ] = 3'd0;
    assign memory1b[163 ] = 3'd2;
    assign memory1b[164 ] = 3'd0;
    assign memory1b[165 ] = 3'd0;
    assign memory1b[166 ] = 3'd0;
    assign memory1b[167 ] = 3'd0;
    assign memory1b[168 ] = 3'd1;
    assign memory1b[169 ] = 3'd2;
    assign memory1b[170 ] = 3'd4;
    assign memory1b[171 ] = 3'd0;
    assign memory1b[172 ] = 3'd2;
    assign memory1b[173 ] = 3'd2;
    assign memory1b[174 ] = 3'd0;
    assign memory1b[175 ] = 3'd0;
    assign memory1b[176 ] = 3'd4;
    assign memory1b[177 ] = 3'd0;
    assign memory1b[178 ] = 3'd0;
    assign memory1b[179 ] = 3'd0;
    assign memory1b[180 ] = 3'd3;
    assign memory1b[181 ] = 3'd0;
    assign memory1b[182 ] = 3'd0;
    assign memory1b[183 ] = 3'd0;
    assign memory1b[184 ] = 3'd2;
    assign memory1b[185 ] = 3'd2;
    assign memory1b[186 ] = 3'd0;
    assign memory1b[187 ] = 3'd0;
    assign memory1b[188 ] = 3'd0;
    assign memory1b[189 ] = 3'd2;
    assign memory1b[190 ] = 3'd2;
    assign memory1b[191 ] = 3'd4;
    assign memory1b[192 ] = 3'd0;
    assign memory1b[193 ] = 3'd4;
    assign memory1b[194 ] = 3'd2;
    assign memory1b[195 ] = 3'd0;
    assign memory1b[196 ] = 3'd0;
    assign memory1b[197 ] = 3'd0;
    assign memory1b[198 ] = 3'd0;
    assign memory1b[199 ] = 3'd1;
    assign memory1b[200 ] = 3'd2;
    assign memory1b[201 ] = 3'd4;
    assign memory1b[202 ] = 3'd2;
    assign memory1b[203 ] = 3'd2;
    assign memory1b[204 ] = 3'd4;
    assign memory1b[205 ] = 3'd2;
    assign memory1b[206 ] = 3'd1;
    assign memory1b[207 ] = 3'd0;
    assign memory1b[208 ] = 3'd4;
    assign memory1b[209 ] = 3'd3;
    assign memory1b[210 ] = 3'd0;
    assign memory1b[211 ] = 3'd0;
    assign memory1b[212 ] = 3'd2;
    assign memory1b[213 ] = 3'd0;
    assign memory1b[214 ] = 3'd2;
    assign memory1b[215 ] = 3'd0;
    assign memory1b[216 ] = 3'd2;
    assign memory1b[217 ] = 3'd0;
    assign memory1b[218 ] = 3'd2;
    assign memory1b[219 ] = 3'd0;
    assign memory1b[220 ] = 3'd4;
    assign memory1b[221 ] = 3'd0;
    assign memory1b[222 ] = 3'd0;
    assign memory1b[223 ] = 3'd0;
    assign memory1b[224 ] = 3'd2;
    assign memory1b[225 ] = 3'd0;
    assign memory1b[226 ] = 3'd0;
    assign memory1b[227 ] = 3'd2;
    assign memory1b[228 ] = 3'd0;
    assign memory1b[229 ] = 3'd0;
    assign memory1b[230 ] = 3'd0;
    assign memory1b[231 ] = 3'd0;
    assign memory1b[232 ] = 3'd0;
    assign memory1b[233 ] = 3'd4;
    assign memory1b[234 ] = 3'd2;
    assign memory1b[235 ] = 3'd0;
    assign memory1b[236 ] = 3'd4;
    assign memory1b[237 ] = 3'd0;
    assign memory1b[238 ] = 3'd0;
    assign memory1b[239 ] = 3'd2;
    assign memory1b[240 ] = 3'd0;
    assign memory1b[241 ] = 3'd4;
    assign memory1b[242 ] = 3'd4;
    assign memory1b[243 ] = 3'd2;
    assign memory1b[244 ] = 3'd4;
    assign memory1b[245 ] = 3'd3;
    assign memory1b[246 ] = 3'd4;
    assign memory1b[247 ] = 3'd4;
    assign memory1b[248 ] = 3'd2;
    assign memory1b[249 ] = 3'd0;
    assign memory1b[250 ] = 3'd4;
    assign memory1b[251 ] = 3'd0;
    assign memory1b[252 ] = 3'd0;
    assign memory1b[253 ] = 3'd0;
    assign memory1b[254 ] = 3'd0;
    assign memory1b[255 ] = 3'd0;
    assign memory1b[256 ] = 3'd0;
    assign memory1b[257 ] = 3'd2;
    assign memory1b[258 ] = 3'd0;
    assign memory1b[259 ] = 3'd2;
    assign memory1b[260 ] = 3'd4;
    assign memory1b[261 ] = 3'd2;
    assign memory1b[262 ] = 3'd2;
    assign memory1b[263 ] = 3'd0;
    assign memory1b[264 ] = 3'd2;
    assign memory1b[265 ] = 3'd2;
    assign memory1b[266 ] = 3'd3;
    assign memory1b[267 ] = 3'd2;
    assign memory1b[268 ] = 3'd0;
    assign memory1b[269 ] = 3'd0;
    assign memory1b[270 ] = 3'd2;
    assign memory1b[271 ] = 3'd4;
    assign memory1b[272 ] = 3'd4;
    assign memory1b[273 ] = 3'd0;
    assign memory1b[274 ] = 3'd0;
    assign memory1b[275 ] = 3'd4;
    assign memory1b[276 ] = 3'd0;
    assign memory1b[277 ] = 3'd4;
    assign memory1b[278 ] = 3'd4;
    assign memory1b[279 ] = 3'd0;
    assign memory1b[280 ] = 3'd4;
    assign memory1b[281 ] = 3'd4;
    assign memory1b[282 ] = 3'd0;
    assign memory1b[283 ] = 3'd0;
    assign memory1b[284 ] = 3'd1;
    assign memory1b[285 ] = 3'd0;
    assign memory1b[286 ] = 3'd0;
    assign memory1b[287 ] = 3'd0;
    assign memory1b[288 ] = 3'd0;
    assign memory1b[289 ] = 3'd2;
    assign memory1b[290 ] = 3'd4;
    assign memory1b[291 ] = 3'd0;
    assign memory1b[292 ] = 3'd2;
    assign memory1b[293 ] = 3'd2;
    assign memory1b[294 ] = 3'd1;
    assign memory1b[295 ] = 3'd0;
    assign memory1b[296 ] = 3'd1;
    assign memory1b[297 ] = 3'd4;
    assign memory1b[298 ] = 3'd0;
    assign memory1b[299 ] = 3'd4;
    assign memory1b[300 ] = 3'd2;
    assign memory1b[301 ] = 3'd0;
    assign memory1b[302 ] = 3'd2;
    assign memory1b[303 ] = 3'd2;
    assign memory1b[304 ] = 3'd0;
    assign memory1b[305 ] = 3'd4;
    assign memory1b[306 ] = 3'd4;
    assign memory1b[307 ] = 3'd0;
    assign memory1b[308 ] = 3'd0;
    assign memory1b[309 ] = 3'd2;
    assign memory1b[310 ] = 3'd0;
    assign memory1b[311 ] = 3'd0;
    assign memory1b[312 ] = 3'd2;
    assign memory1b[313 ] = 3'd3;
    assign memory1b[314 ] = 3'd0;
    assign memory1b[315 ] = 3'd2;
    assign memory1b[316 ] = 3'd0;
    assign memory1b[317 ] = 3'd2;
    assign memory1b[318 ] = 3'd0;
    assign memory1b[319 ] = 3'd0;
    assign memory1b[320 ] = 3'd4;
    assign memory1b[321 ] = 3'd0;
    assign memory1b[322 ] = 3'd2;
    assign memory1b[323 ] = 3'd2;
    assign memory1b[324 ] = 3'd2;
    assign memory1b[325 ] = 3'd0;
    assign memory1b[326 ] = 3'd0;
    assign memory1b[327 ] = 3'd2;
    assign memory1b[328 ] = 3'd0;
    assign memory1b[329 ] = 3'd1;
    assign memory1b[330 ] = 3'd2;
    assign memory1b[331 ] = 3'd2;
    assign memory1b[332 ] = 3'd0;
    assign memory1b[333 ] = 3'd2;
    assign memory1b[334 ] = 3'd0;
    assign memory1b[335 ] = 3'd2;
    assign memory1b[336 ] = 3'd4;
    assign memory1b[337 ] = 3'd2;
    assign memory1b[338 ] = 3'd0;
    assign memory1b[339 ] = 3'd2;
    assign memory1b[340 ] = 3'd0;
    assign memory1b[341 ] = 3'd2;
    assign memory1b[342 ] = 3'd2;
    assign memory1b[343 ] = 3'd2;
    assign memory1b[344 ] = 3'd0;
    assign memory1b[345 ] = 3'd0;
    assign memory1b[346 ] = 3'd0;
    assign memory1b[347 ] = 3'd0;
    assign memory1b[348 ] = 3'd0;
    assign memory1b[349 ] = 3'd2;
    assign memory1b[350 ] = 3'd0;
    assign memory1b[351 ] = 3'd4;
    assign memory1b[352 ] = 3'd2;
    assign memory1b[353 ] = 3'd2;
    assign memory1b[354 ] = 3'd0;
    assign memory1b[355 ] = 3'd2;
    assign memory1b[356 ] = 3'd4;
    assign memory1b[357 ] = 3'd2;
    assign memory1b[358 ] = 3'd0;
    assign memory1b[359 ] = 3'd2;
    assign memory1b[360 ] = 3'd2;
    assign memory1b[361 ] = 3'd0;
    assign memory1b[362 ] = 3'd4;
    assign memory1b[363 ] = 3'd0;
    assign memory1b[364 ] = 3'd4;
    assign memory1b[365 ] = 3'd0;
    assign memory1b[366 ] = 3'd4;
    assign memory1b[367 ] = 3'd2;
    assign memory1b[368 ] = 3'd1;
    assign memory1b[369 ] = 3'd4;
    assign memory1b[370 ] = 3'd0;
    assign memory1b[371 ] = 3'd2;
    assign memory1b[372 ] = 3'd0;
    assign memory1b[373 ] = 3'd1;
    assign memory1b[374 ] = 3'd4;
    assign memory1b[375 ] = 3'd2;
    assign memory1b[376 ] = 3'd0;
    assign memory1b[377 ] = 3'd2;
    assign memory1b[378 ] = 3'd1;
    assign memory1b[379 ] = 3'd0;
    assign memory1b[380 ] = 3'd2;
    assign memory1b[381 ] = 3'd2;
    assign memory1b[382 ] = 3'd3;
    assign memory1b[383 ] = 3'd4;
    assign memory1b[384 ] = 3'd0;
    assign memory1b[385 ] = 3'd4;
    assign memory1b[386 ] = 3'd2;
    assign memory1b[387 ] = 3'd2;
    assign memory1b[388 ] = 3'd0;
    assign memory1b[389 ] = 3'd0;
    assign memory1b[390 ] = 3'd2;
    assign memory1b[391 ] = 3'd2;
    assign memory1b[392 ] = 3'd0;
    assign memory1b[393 ] = 3'd0;
    assign memory1b[394 ] = 3'd1;
    assign memory1b[395 ] = 3'd2;
    assign memory1b[396 ] = 3'd2;
    assign memory1b[397 ] = 3'd2;
    assign memory1b[398 ] = 3'd3;
    assign memory1b[399 ] = 3'd4;
    assign memory1b[400 ] = 3'd2;
    assign memory1b[401 ] = 3'd4;
    assign memory1b[402 ] = 3'd2;
    assign memory1b[403 ] = 3'd2;
    assign memory1b[404 ] = 3'd4;
    assign memory1b[405 ] = 3'd0;
    assign memory1b[406 ] = 3'd0;
    assign memory1b[407 ] = 3'd4;
    assign memory1b[408 ] = 3'd4;
    assign memory1b[409 ] = 3'd0;
    assign memory1b[410 ] = 3'd4;
    assign memory1b[411 ] = 3'd0;
    assign memory1b[412 ] = 3'd0;
    assign memory1b[413 ] = 3'd0;
    assign memory1b[414 ] = 3'd0;
    assign memory1b[415 ] = 3'd0;
    assign memory1b[416 ] = 3'd0;
    assign memory1b[417 ] = 3'd2;
    assign memory1b[418 ] = 3'd0;
    assign memory1b[419 ] = 3'd0;
    assign memory1b[420 ] = 3'd0;
    assign memory1b[421 ] = 3'd0;
    assign memory1b[422 ] = 3'd0;
    assign memory1b[423 ] = 3'd0;
    assign memory1b[424 ] = 3'd0;
    assign memory1b[425 ] = 3'd0;
    assign memory1b[426 ] = 3'd2;
    assign memory1b[427 ] = 3'd0;
    assign memory1b[428 ] = 3'd4;
    assign memory1b[429 ] = 3'd2;
    assign memory1b[430 ] = 3'd0;
    assign memory1b[431 ] = 3'd2;
    assign memory1b[432 ] = 3'd0;
    assign memory1b[433 ] = 3'd0;
    assign memory1b[434 ] = 3'd0;
    assign memory1b[435 ] = 3'd0;
    assign memory1b[436 ] = 3'd2;
    assign memory1b[437 ] = 3'd2;
    assign memory1b[438 ] = 3'd0;
    assign memory1b[439 ] = 3'd0;
    assign memory1b[440 ] = 3'd0;
    assign memory1b[441 ] = 3'd0;
    assign memory1b[442 ] = 3'd0;
    assign memory1b[443 ] = 3'd0;
    assign memory1b[444 ] = 3'd2;
    assign memory1b[445 ] = 3'd2;
    assign memory1b[446 ] = 3'd4;
    assign memory1b[447 ] = 3'd0;
    assign memory1b[448 ] = 3'd0;
    assign memory1b[449 ] = 3'd0;
    assign memory1b[450 ] = 3'd1;
    assign memory1b[451 ] = 3'd4;
    assign memory1b[452 ] = 3'd2;
    assign memory1b[453 ] = 3'd3;
    assign memory1b[454 ] = 3'd0;
    assign memory1b[455 ] = 3'd0;
    assign memory1b[456 ] = 3'd0;
    assign memory1b[457 ] = 3'd0;
    assign memory1b[458 ] = 3'd0;
    assign memory1b[459 ] = 3'd0;
    assign memory1b[460 ] = 3'd0;
    assign memory1b[461 ] = 3'd4;
    assign memory1b[462 ] = 3'd2;
    assign memory1b[463 ] = 3'd0;
    assign memory1b[464 ] = 3'd0;
    assign memory1b[465 ] = 3'd0;
    assign memory1b[466 ] = 3'd0;
    assign memory1b[467 ] = 3'd1;
    assign memory1b[468 ] = 3'd2;
    assign memory1b[469 ] = 3'd4;
    assign memory1b[470 ] = 3'd2;
    assign memory1b[471 ] = 3'd2;
    assign memory1b[472 ] = 3'd4;
    assign memory1b[473 ] = 3'd2;
    assign memory1b[474 ] = 3'd1;
    assign memory1b[475 ] = 3'd0;
    assign memory1b[476 ] = 3'd4;
    assign memory1b[477 ] = 3'd3;
    assign memory1b[478 ] = 3'd0;
    assign memory1b[479 ] = 3'd0;
    assign memory1b[480 ] = 3'd3;
    assign memory1b[481 ] = 3'd0;
    assign memory1b[482 ] = 3'd2;
    assign memory1b[483 ] = 3'd0;
    assign memory1b[484 ] = 3'd2;
    assign memory1b[485 ] = 3'd0;
    assign memory1b[486 ] = 3'd0;
    assign memory1b[487 ] = 3'd0;
    assign memory1b[488 ] = 3'd2;
    assign memory1b[489 ] = 3'd0;
    assign memory1b[490 ] = 3'd0;
    assign memory1b[491 ] = 3'd0;
    assign memory1b[492 ] = 3'd0;
    assign memory1b[493 ] = 3'd2;
    assign memory1b[494 ] = 3'd1;
    assign memory1b[495 ] = 3'd0;
    assign memory1b[496 ] = 3'd2;
    assign memory1b[497 ] = 3'd0;
    assign memory1b[498 ] = 3'd0;
    assign memory1b[499 ] = 3'd0;
    assign memory1b[500 ] = 3'd2;
    assign memory1b[501 ] = 3'd0;
    assign memory1b[502 ] = 3'd2;
    assign memory1b[503 ] = 3'd0;
    assign memory1b[504 ] = 3'd2;
    assign memory1b[505 ] = 3'd3;
    assign memory1b[506 ] = 3'd2;
    assign memory1b[507 ] = 3'd2;
    assign memory1b[508 ] = 3'd2;
    assign memory1b[509 ] = 3'd0;
    assign memory1b[510 ] = 3'd0;
    assign memory1b[511 ] = 3'd0;
    assign memory1b[512 ] = 3'd0;
    assign memory1b[513 ] = 3'd0;
    assign memory1b[514 ] = 3'd0;
    assign memory1b[515 ] = 3'd0;
    assign memory1b[516 ] = 3'd0;
    assign memory1b[517 ] = 3'd0;
    assign memory1b[518 ] = 3'd0;
    assign memory1b[519 ] = 3'd0;
    assign memory1b[520 ] = 3'd2;
    assign memory1b[521 ] = 3'd2;
    assign memory1b[522 ] = 3'd0;
    assign memory1b[523 ] = 3'd2;
    assign memory1b[524 ] = 3'd2;
    assign memory1b[525 ] = 3'd0;
    assign memory1b[526 ] = 3'd0;
    assign memory1b[527 ] = 3'd0;
    assign memory1b[528 ] = 3'd0;
    assign memory1b[529 ] = 3'd0;
    assign memory1b[530 ] = 3'd2;
    assign memory1b[531 ] = 3'd0;
    assign memory1b[532 ] = 3'd0;
    assign memory1b[533 ] = 3'd0;
    assign memory1b[534 ] = 3'd0;
    assign memory1b[535 ] = 3'd2;
    assign memory1b[536 ] = 3'd0;
    assign memory1b[537 ] = 3'd0;
    assign memory1b[538 ] = 3'd0;
    assign memory1b[539 ] = 3'd0;
    assign memory1b[540 ] = 3'd0;
    assign memory1b[541 ] = 3'd2;
    assign memory1b[542 ] = 3'd0;
    assign memory1b[543 ] = 3'd3;
    assign memory1b[544 ] = 3'd2;
    assign memory1b[545 ] = 3'd2;
    assign memory1b[546 ] = 3'd0;
    assign memory1b[547 ] = 3'd4;
    assign memory1b[548 ] = 3'd4;
    assign memory1b[549 ] = 3'd2;
    assign memory1b[550 ] = 3'd0;
    assign memory1b[551 ] = 3'd0;
    assign memory1b[552 ] = 3'd1;
    assign memory1b[553 ] = 3'd0;
    assign memory1b[554 ] = 3'd4;
    assign memory1b[555 ] = 3'd0;
    assign memory1b[556 ] = 3'd2;
    assign memory1b[557 ] = 3'd2;
    assign memory1b[558 ] = 3'd0;
    assign memory1b[559 ] = 3'd0;
    assign memory1b[560 ] = 3'd0;
    assign memory1b[561 ] = 3'd1;
    assign memory1b[562 ] = 3'd0;
    assign memory1b[563 ] = 3'd0;
    assign memory1b[564 ] = 3'd0;
    assign memory1b[565 ] = 3'd0;
    assign memory1b[566 ] = 3'd0;
    assign memory1b[567 ] = 3'd0;
    assign memory1b[568 ] = 3'd0;
    assign memory1b[569 ] = 3'd4;
    assign memory1b[570 ] = 3'd4;
    assign memory1b[571 ] = 3'd0;
    assign memory1b[572 ] = 3'd2;
    assign memory1b[573 ] = 3'd0;
    assign memory1b[574 ] = 3'd0;
    assign memory1b[575 ] = 3'd0;
    assign memory1b[576 ] = 3'd4;
    assign memory1b[577 ] = 3'd0;
    assign memory1b[578 ] = 3'd4;
    assign memory1b[579 ] = 3'd2;
    assign memory1b[580 ] = 3'd4;
    assign memory1b[581 ] = 3'd2;
    assign memory1b[582 ] = 3'd0;
    assign memory1b[583 ] = 3'd0;
    assign memory1b[584 ] = 3'd0;
    assign memory1b[585 ] = 3'd0;
    assign memory1b[586 ] = 3'd0;
    assign memory1b[587 ] = 3'd2;
    assign memory1b[588 ] = 3'd0;
    assign memory1b[589 ] = 3'd4;
    assign memory1b[590 ] = 3'd4;
    assign memory1b[591 ] = 3'd4;
    assign memory1b[592 ] = 3'd0;
    assign memory1b[593 ] = 3'd4;
    assign memory1b[594 ] = 3'd0;
    assign memory1b[595 ] = 3'd4;
    assign memory1b[596 ] = 3'd2;
    assign memory1b[597 ] = 3'd0;
    assign memory1b[598 ] = 3'd0;
    assign memory1b[599 ] = 3'd0;
    assign memory1b[600 ] = 3'd2;
    assign memory1b[601 ] = 3'd4;
    assign memory1b[602 ] = 3'd0;
    assign memory1b[603 ] = 3'd2;
    assign memory1b[604 ] = 3'd2;
    assign memory1b[605 ] = 3'd0;
    assign memory1b[606 ] = 3'd0;
    assign memory1b[607 ] = 3'd4;
    assign memory1b[608 ] = 3'd4;
    assign memory1b[609 ] = 3'd0;
    assign memory1b[610 ] = 3'd2;
    assign memory1b[611 ] = 3'd0;
    assign memory1b[612 ] = 3'd4;
    assign memory1b[613 ] = 3'd4;
    assign memory1b[614 ] = 3'd0;
    assign memory1b[615 ] = 3'd0;
    assign memory1b[616 ] = 3'd0;
    assign memory1b[617 ] = 3'd2;
    assign memory1b[618 ] = 3'd2;
    assign memory1b[619 ] = 3'd0;
    assign memory1b[620 ] = 3'd2;
    assign memory1b[621 ] = 3'd1;
    assign memory1b[622 ] = 3'd1;
    assign memory1b[623 ] = 3'd2;
    assign memory1b[624 ] = 3'd0;
    assign memory1b[625 ] = 3'd0;
    assign memory1b[626 ] = 3'd0;
    assign memory1b[627 ] = 3'd0;
    assign memory1b[628 ] = 3'd0;
    assign memory1b[629 ] = 3'd0;
    assign memory1b[630 ] = 3'd0;
    assign memory1b[631 ] = 3'd0;
    assign memory1b[632 ] = 3'd2;
    assign memory1b[633 ] = 3'd2;
    assign memory1b[634 ] = 3'd1;
    assign memory1b[635 ] = 3'd0;
    assign memory1b[636 ] = 3'd0;
    assign memory1b[637 ] = 3'd0;
    assign memory1b[638 ] = 3'd0;
    assign memory1b[639 ] = 3'd2;
    assign memory1b[640 ] = 3'd3;
    assign memory1b[641 ] = 3'd4;
    assign memory1b[642 ] = 3'd0;
    assign memory1b[643 ] = 3'd2;
    assign memory1b[644 ] = 3'd0;
    assign memory1b[645 ] = 3'd0;
    assign memory1b[646 ] = 3'd0;
    assign memory1b[647 ] = 3'd1;
    assign memory1b[648 ] = 3'd0;
    assign memory1b[649 ] = 3'd0;
    assign memory1b[650 ] = 3'd0;
    assign memory1b[651 ] = 3'd0;
    assign memory1b[652 ] = 3'd0;
    assign memory1b[653 ] = 3'd2;
    assign memory1b[654 ] = 3'd0;
    assign memory1b[655 ] = 3'd0;
    assign memory1b[656 ] = 3'd0;
    assign memory1b[657 ] = 3'd4;
    assign memory1b[658 ] = 3'd0;
    assign memory1b[659 ] = 3'd0;
    assign memory1b[660 ] = 3'd1;
    assign memory1b[661 ] = 3'd4;
    assign memory1b[662 ] = 3'd0;
    assign memory1b[663 ] = 3'd0;
    assign memory1b[664 ] = 3'd2;
    assign memory1b[665 ] = 3'd0;
    assign memory1b[666 ] = 3'd0;
    assign memory1b[667 ] = 3'd4;
    assign memory1b[668 ] = 3'd0;
    assign memory1b[669 ] = 3'd0;
    assign memory1b[670 ] = 3'd2;
    assign memory1b[671 ] = 3'd2;
    assign memory1b[672 ] = 3'd4;
    assign memory1b[673 ] = 3'd4;
    assign memory1b[674 ] = 3'd0;
    assign memory1b[675 ] = 3'd4;
    assign memory1b[676 ] = 3'd0;
    assign memory1b[677 ] = 3'd2;
    assign memory1b[678 ] = 3'd1;
    assign memory1b[679 ] = 3'd4;
    assign memory1b[680 ] = 3'd2;
    assign memory1b[681 ] = 3'd2;
    assign memory1b[682 ] = 3'd4;
    assign memory1b[683 ] = 3'd0;
    assign memory1b[684 ] = 3'd0;
    assign memory1b[685 ] = 3'd4;
    assign memory1b[686 ] = 3'd0;
    assign memory1b[687 ] = 3'd0;
    assign memory1b[688 ] = 3'd0;
    assign memory1b[689 ] = 3'd1;
    assign memory1b[690 ] = 3'd0;
    assign memory1b[691 ] = 3'd0;
    assign memory1b[692 ] = 3'd0;
    assign memory1b[693 ] = 3'd0;
    assign memory1b[694 ] = 3'd2;
    assign memory1b[695 ] = 3'd4;
    assign memory1b[696 ] = 3'd0;
    assign memory1b[697 ] = 3'd2;
    assign memory1b[698 ] = 3'd0;
    assign memory1b[699 ] = 3'd2;
    assign memory1b[700 ] = 3'd4;
    assign memory1b[701 ] = 3'd0;
    assign memory1b[702 ] = 3'd2;
    assign memory1b[703 ] = 3'd2;
    assign memory1b[704 ] = 3'd0;
    assign memory1b[705 ] = 3'd0;
    assign memory1b[706 ] = 3'd4;
    assign memory1b[707 ] = 3'd0;
    assign memory1b[708 ] = 3'd4;
    assign memory1b[709 ] = 3'd2;
    assign memory1b[710 ] = 3'd4;
    assign memory1b[711 ] = 3'd2;
    assign memory1b[712 ] = 3'd0;
    assign memory1b[713 ] = 3'd0;
    assign memory1b[714 ] = 3'd0;
    assign memory1b[715 ] = 3'd0;
    assign memory1b[716 ] = 3'd0;
    assign memory1b[717 ] = 3'd2;
    assign memory1b[718 ] = 3'd0;
    assign memory1b[719 ] = 3'd4;
    assign memory1b[720 ] = 3'd4;
    assign memory1b[721 ] = 3'd4;
    assign memory1b[722 ] = 3'd0;
    assign memory1b[723 ] = 3'd4;
    assign memory1b[724 ] = 3'd0;
    assign memory1b[725 ] = 3'd4;
    assign memory1b[726 ] = 3'd2;
    assign memory1b[727 ] = 3'd0;
    assign memory1b[728 ] = 3'd0;
    assign memory1b[729 ] = 3'd0;
    assign memory1b[730 ] = 3'd2;
    assign memory1b[731 ] = 3'd4;
    assign memory1b[732 ] = 3'd0;
    assign memory1b[733 ] = 3'd2;
    assign memory1b[734 ] = 3'd2;
    assign memory1b[735 ] = 3'd0;
    assign memory1b[736 ] = 3'd0;
    assign memory1b[737 ] = 3'd0;
    assign memory1b[738 ] = 3'd0;
    assign memory1b[739 ] = 3'd0;
    assign memory1b[740 ] = 3'd0;
    assign memory1b[741 ] = 3'd1;
    assign memory1b[742 ] = 3'd0;
    assign memory1b[743 ] = 3'd0;
    assign memory1b[744 ] = 3'd0;
    assign memory1b[745 ] = 3'd0;
    assign memory1b[746 ] = 3'd4;
    assign memory1b[747 ] = 3'd2;
    assign memory1b[748 ] = 3'd1;
    assign memory1b[749 ] = 3'd2;
    assign memory1b[750 ] = 3'd0;
    assign memory1b[751 ] = 3'd4;
    assign memory1b[752 ] = 3'd0;
    assign memory1b[753 ] = 3'd1;
    assign memory1b[754 ] = 3'd4;
    assign memory1b[755 ] = 3'd0;
    assign memory1b[756 ] = 3'd0;
    assign memory1b[757 ] = 3'd0;
    assign memory1b[758 ] = 3'd0;
    assign memory1b[759 ] = 3'd4;
    assign memory1b[760 ] = 3'd0;
    assign memory1b[761 ] = 3'd2;
    assign memory1b[762 ] = 3'd2;
    assign memory1b[763 ] = 3'd2;
    assign memory1b[764 ] = 3'd1;
    assign memory1b[765 ] = 3'd4;
    assign memory1b[766 ] = 3'd0;
    assign memory1b[767 ] = 3'd2;
    assign memory1b[768 ] = 3'd2;
    assign memory1b[769 ] = 3'd0;
    assign memory1b[770 ] = 3'd2;
    assign memory1b[771 ] = 3'd2;
    assign memory1b[772 ] = 3'd0;
    assign memory1b[773 ] = 3'd2;
    assign memory1b[774 ] = 3'd0;
    assign memory1b[775 ] = 3'd2;
    assign memory1b[776 ] = 3'd0;
    assign memory1b[777 ] = 3'd4;
    assign memory1b[778 ] = 3'd2;
    assign memory1b[779 ] = 3'd0;
    assign memory1b[780 ] = 3'd1;
    assign memory1b[781 ] = 3'd0;
    assign memory1b[782 ] = 3'd2;
    assign memory1b[783 ] = 3'd3;
    assign memory1b[784 ] = 3'd0;
    assign memory1b[785 ] = 3'd4;
    assign memory1b[786 ] = 3'd4;
    assign memory1b[787 ] = 3'd2;
    assign memory1b[788 ] = 3'd0;
    assign memory1b[789 ] = 3'd2;
    assign memory1b[790 ] = 3'd0;
    assign memory1b[791 ] = 3'd2;
    assign memory1b[792 ] = 3'd0;
    assign memory1b[793 ] = 3'd0;
    assign memory1b[794 ] = 3'd4;
    assign memory1b[795 ] = 3'd2;
    assign memory1b[796 ] = 3'd2;
    assign memory1b[797 ] = 3'd0;
    assign memory1b[798 ] = 3'd2;
    assign memory1b[799 ] = 3'd4;
    assign memory1b[800 ] = 3'd2;
    assign memory1b[801 ] = 3'd2;
    assign memory1b[802 ] = 3'd0;
    assign memory1b[803 ] = 3'd0;
    assign memory1b[804 ] = 3'd1;
    assign memory1b[805 ] = 3'd0;
    assign memory1b[806 ] = 3'd0;
    assign memory1b[807 ] = 3'd0;
    assign memory1b[808 ] = 3'd2;
    assign memory1b[809 ] = 3'd2;
    assign memory1b[810 ] = 3'd0;
    assign memory1b[811 ] = 3'd2;
    assign memory1b[812 ] = 3'd2;
    assign memory1b[813 ] = 3'd0;
    assign memory1b[814 ] = 3'd2;
    assign memory1b[815 ] = 3'd0;
    assign memory1b[816 ] = 3'd2;
    assign memory1b[817 ] = 3'd0;
    assign memory1b[818 ] = 3'd0;
    assign memory1b[819 ] = 3'd2;
    assign memory1b[820 ] = 3'd0;
    assign memory1b[821 ] = 3'd4;
    assign memory1b[822 ] = 3'd2;
    assign memory1b[823 ] = 3'd0;
    assign memory1b[824 ] = 3'd0;
    assign memory1b[825 ] = 3'd0;
    assign memory1b[826 ] = 3'd0;
    assign memory1b[827 ] = 3'd0;
    assign memory1b[828 ] = 3'd2;
    assign memory1b[829 ] = 3'd2;
    assign memory1b[830 ] = 3'd0;
    assign memory1b[831 ] = 3'd4;
    assign memory1b[832 ] = 3'd0;
    assign memory1b[833 ] = 3'd0;
    assign memory1b[834 ] = 3'd0;
    assign memory1b[835 ] = 3'd0;
    assign memory1b[836 ] = 3'd0;
    assign memory1b[837 ] = 3'd0;
    assign memory1b[838 ] = 3'd0;
    assign memory1b[839 ] = 3'd0;
    assign memory1b[840 ] = 3'd0;
    assign memory1b[841 ] = 3'd1;
    assign memory1b[842 ] = 3'd1;
    assign memory1b[843 ] = 3'd0;
    assign memory1b[844 ] = 3'd2;
    assign memory1b[845 ] = 3'd0;
    assign memory1b[846 ] = 3'd0;
    assign memory1b[847 ] = 3'd0;
    assign memory1b[848 ] = 3'd0;
    assign memory1b[849 ] = 3'd0;
    assign memory1b[850 ] = 3'd4;
    assign memory1b[851 ] = 3'd0;
    assign memory1b[852 ] = 3'd0;
    assign memory1b[853 ] = 3'd0;
    assign memory1b[854 ] = 3'd0;
    assign memory1b[855 ] = 3'd4;
    assign memory1b[856 ] = 3'd2;
    assign memory1b[857 ] = 3'd0;
    assign memory1b[858 ] = 3'd3;
    assign memory1b[859 ] = 3'd2;
    assign memory1b[860 ] = 3'd0;
    assign memory1b[861 ] = 3'd0;
    assign memory1b[862 ] = 3'd0;
    assign memory1b[863 ] = 3'd1;
    assign memory1b[864 ] = 3'd4;
    assign memory1b[865 ] = 3'd4;
    assign memory1b[866 ] = 3'd0;
    assign memory1b[867 ] = 3'd2;
    assign memory1b[868 ] = 3'd0;
    assign memory1b[869 ] = 3'd0;
    assign memory1b[870 ] = 3'd0;
    assign memory1b[871 ] = 3'd2;
    assign memory1b[872 ] = 3'd0;
    assign memory1b[873 ] = 3'd0;
    assign memory1b[874 ] = 3'd3;
    assign memory1b[875 ] = 3'd2;
    assign memory1b[876 ] = 3'd2;
    assign memory1b[877 ] = 3'd4;
    assign memory1b[878 ] = 3'd2;
    assign memory1b[879 ] = 3'd4;
    assign memory1b[880 ] = 3'd0;
    assign memory1b[881 ] = 3'd4;
    assign memory1b[882 ] = 3'd2;
    assign memory1b[883 ] = 3'd0;
    assign memory1b[884 ] = 3'd0;
    assign memory1b[885 ] = 3'd0;
    assign memory1b[886 ] = 3'd1;
    assign memory1b[887 ] = 3'd0;
    assign memory1b[888 ] = 3'd4;
    assign memory1b[889 ] = 3'd0;
    assign memory1b[890 ] = 3'd2;
    assign memory1b[891 ] = 3'd0;
    assign memory1b[892 ] = 3'd2;
    assign memory1b[893 ] = 3'd0;
    assign memory1b[894 ] = 3'd0;
    assign memory1b[895 ] = 3'd0;
    assign memory1b[896 ] = 3'd2;
    assign memory1b[897 ] = 3'd4;
    assign memory1b[898 ] = 3'd0;
    assign memory1b[899 ] = 3'd2;
    assign memory1b[900 ] = 3'd1;
    assign memory1b[901 ] = 3'd0;
    assign memory1b[902 ] = 3'd1;
    assign memory1b[903 ] = 3'd0;
    assign memory1b[904 ] = 3'd0;
    assign memory1b[905 ] = 3'd0;
    assign memory1b[906 ] = 3'd2;
    assign memory1b[907 ] = 3'd4;
    assign memory1b[908 ] = 3'd2;
    assign memory1b[909 ] = 3'd0;
    assign memory1b[910 ] = 3'd0;
    assign memory1b[911 ] = 3'd4;
    assign memory1b[912 ] = 3'd0;
    assign memory1b[913 ] = 3'd2;
    assign memory1b[914 ] = 3'd0;
    assign memory1b[915 ] = 3'd2;
    assign memory1b[916 ] = 3'd0;
    assign memory1b[917 ] = 3'd2;
    assign memory1b[918 ] = 3'd2;
    assign memory1b[919 ] = 3'd4;
    assign memory1b[920 ] = 3'd0;
    assign memory1b[921 ] = 3'd3;
    assign memory1b[922 ] = 3'd4;
    assign memory1b[923 ] = 3'd0;
    assign memory1b[924 ] = 3'd0;
    assign memory1b[925 ] = 3'd0;
    assign memory1b[926 ] = 3'd2;
    assign memory1b[927 ] = 3'd0;
    assign memory1b[928 ] = 3'd0;
    assign memory1b[929 ] = 3'd0;
    assign memory1b[930 ] = 3'd2;
    assign memory1b[931 ] = 3'd2;
    assign memory1b[932 ] = 3'd0;
    assign memory1b[933 ] = 3'd2;
    assign memory1b[934 ] = 3'd2;
    assign memory1b[935 ] = 3'd0;
    assign memory1b[936 ] = 3'd0;
    assign memory1b[937 ] = 3'd0;
    assign memory1b[938 ] = 3'd0;
    assign memory1b[939 ] = 3'd0;
    assign memory1b[940 ] = 3'd2;
    assign memory1b[941 ] = 3'd0;
    assign memory1b[942 ] = 3'd0;
    assign memory1b[943 ] = 3'd0;
    assign memory1b[944 ] = 3'd0;
    assign memory1b[945 ] = 3'd2;
    assign memory1b[946 ] = 3'd0;
    assign memory1b[947 ] = 3'd0;
    assign memory1b[948 ] = 3'd0;
    assign memory1b[949 ] = 3'd0;
    assign memory1b[950 ] = 3'd0;
    assign memory1b[951 ] = 3'd2;
    assign memory1b[952 ] = 3'd0;
    assign memory1b[953 ] = 3'd3;
    assign memory1b[954 ] = 3'd0;
    assign memory1b[955 ] = 3'd0;
    assign memory1b[956 ] = 3'd0;
    assign memory1b[957 ] = 3'd0;
    assign memory1b[958 ] = 3'd0;
    assign memory1b[959 ] = 3'd0;
    assign memory1b[960 ] = 3'd0;
    assign memory1b[961 ] = 3'd0;
    assign memory1b[962 ] = 3'd4;
    assign memory1b[963 ] = 3'd4;
    assign memory1b[964 ] = 3'd0;
    assign memory1b[965 ] = 3'd4;
    assign memory1b[966 ] = 3'd0;
    assign memory1b[967 ] = 3'd0;
    assign memory1b[968 ] = 3'd0;
    assign memory1b[969 ] = 3'd2;
    assign memory1b[970 ] = 3'd2;
    assign memory1b[971 ] = 3'd0;
    assign memory1b[972 ] = 3'd0;
    assign memory1b[973 ] = 3'd1;
    assign memory1b[974 ] = 3'd1;
    assign memory1b[975 ] = 3'd0;
    assign memory1b[976 ] = 3'd0;
    assign memory1b[977 ] = 3'd0;
    assign memory1b[978 ] = 3'd0;
    assign memory1b[979 ] = 3'd4;
    assign memory1b[980 ] = 3'd2;
    assign memory1b[981 ] = 3'd2;
    assign memory1b[982 ] = 3'd0;
    assign memory1b[983 ] = 3'd0;
    assign memory1b[984 ] = 3'd0;
    assign memory1b[985 ] = 3'd0;
    assign memory1b[986 ] = 3'd0;
    assign memory1b[987 ] = 3'd0;
    assign memory1b[988 ] = 3'd0;
    assign memory1b[989 ] = 3'd0;
    assign memory1b[990 ] = 3'd0;
    assign memory1b[991 ] = 3'd2;
    assign memory1b[992 ] = 3'd2;
    assign memory1b[993 ] = 3'd2;
    assign memory1b[994 ] = 3'd0;
    assign memory1b[995 ] = 3'd0;
    assign memory1b[996 ] = 3'd4;
    assign memory1b[997 ] = 3'd0;
    assign memory1b[998 ] = 3'd2;
    assign memory1b[999 ] = 3'd0;
    assign memory1b[1000] = 3'd2;
    assign memory1b[1001] = 3'd4;
    assign memory1b[1002] = 3'd2;
    assign memory1b[1003] = 3'd2;
    assign memory1b[1004] = 3'd4;
    assign memory1b[1005] = 3'd4;
    assign memory1b[1006] = 3'd0;
    assign memory1b[1007] = 3'd2;
    assign memory1b[1008] = 3'd0;
    assign memory1b[1009] = 3'd0;
    assign memory1b[1010] = 3'd4;
    assign memory1b[1011] = 3'd0;
    assign memory1b[1012] = 3'd2;
    assign memory1b[1013] = 3'd0;
    assign memory1b[1014] = 3'd1;
    assign memory1b[1015] = 3'd3;
    assign memory1b[1016] = 3'd0;
    assign memory1b[1017] = 3'd2;
    assign memory1b[1018] = 3'd0;
    assign memory1b[1019] = 3'd2;
    assign memory1b[1020] = 3'd0;
    assign memory1b[1021] = 3'd0;
    assign memory1b[1022] = 3'd0;
    assign memory1b[1023] = 3'd0;

    assign memory3a[0   ] = 3'd0;
    assign memory3a[1   ] = 3'd1;
    assign memory3a[2   ] = 3'd2;
    assign memory3a[3   ] = 3'd2;
    assign memory3a[4   ] = 3'd1;
    assign memory3a[5   ] = 3'd2;
    assign memory3a[6   ] = 3'd2;
    assign memory3a[7   ] = 3'd2;
    assign memory3a[8   ] = 3'd0;
    assign memory3a[9   ] = 3'd2;
    assign memory3a[10  ] = 3'd0;
    assign memory3a[11  ] = 3'd2;
    assign memory3a[12  ] = 3'd2;
    assign memory3a[13  ] = 3'd1;
    assign memory3a[14  ] = 3'd2;
    assign memory3a[15  ] = 3'd2;
    assign memory3a[16  ] = 3'd2;
    assign memory3a[17  ] = 3'd2;
    assign memory3a[18  ] = 3'd2;
    assign memory3a[19  ] = 3'd0;
    assign memory3a[20  ] = 3'd2;
    assign memory3a[21  ] = 3'd0;
    assign memory3a[22  ] = 3'd2;
    assign memory3a[23  ] = 3'd2;
    assign memory3a[24  ] = 3'd2;
    assign memory3a[25  ] = 3'd2;
    assign memory3a[26  ] = 3'd0;
    assign memory3a[27  ] = 3'd2;
    assign memory3a[28  ] = 3'd2;
    assign memory3a[29  ] = 3'd2;
    assign memory3a[30  ] = 3'd2;
    assign memory3a[31  ] = 3'd2;
    assign memory3a[32  ] = 3'd1;
    assign memory3a[33  ] = 3'd2;
    assign memory3a[34  ] = 3'd2;
    assign memory3a[35  ] = 3'd1;
    assign memory3a[36  ] = 3'd2;
    assign memory3a[37  ] = 3'd2;
    assign memory3a[38  ] = 3'd2;
    assign memory3a[39  ] = 3'd2;
    assign memory3a[40  ] = 3'd0;
    assign memory3a[41  ] = 3'd2;
    assign memory3a[42  ] = 3'd0;
    assign memory3a[43  ] = 3'd1;
    assign memory3a[44  ] = 3'd2;
    assign memory3a[45  ] = 3'd1;
    assign memory3a[46  ] = 3'd2;
    assign memory3a[47  ] = 3'd2;
    assign memory3a[48  ] = 3'd2;
    assign memory3a[49  ] = 3'd2;
    assign memory3a[50  ] = 3'd0;
    assign memory3a[51  ] = 3'd1;
    assign memory3a[52  ] = 3'd2;
    assign memory3a[53  ] = 3'd2;
    assign memory3a[54  ] = 3'd2;
    assign memory3a[55  ] = 3'd2;
    assign memory3a[56  ] = 3'd2;
    assign memory3a[57  ] = 3'd0;
    assign memory3a[58  ] = 3'd1;
    assign memory3a[59  ] = 3'd2;
    assign memory3a[60  ] = 3'd2;
    assign memory3a[61  ] = 3'd0;
    assign memory3a[62  ] = 3'd2;
    assign memory3a[63  ] = 3'd2;
    assign memory3a[64  ] = 3'd0;
    assign memory3a[65  ] = 3'd2;
    assign memory3a[66  ] = 3'd2;
    assign memory3a[67  ] = 3'd1;
    assign memory3a[68  ] = 3'd2;
    assign memory3a[69  ] = 3'd2;
    assign memory3a[70  ] = 3'd0;
    assign memory3a[71  ] = 3'd2;
    assign memory3a[72  ] = 3'd2;
    assign memory3a[73  ] = 3'd2;
    assign memory3a[74  ] = 3'd2;
    assign memory3a[75  ] = 3'd1;
    assign memory3a[76  ] = 3'd2;
    assign memory3a[77  ] = 3'd2;
    assign memory3a[78  ] = 3'd2;
    assign memory3a[79  ] = 3'd2;
    assign memory3a[80  ] = 3'd2;
    assign memory3a[81  ] = 3'd0;
    assign memory3a[82  ] = 3'd2;
    assign memory3a[83  ] = 3'd1;
    assign memory3a[84  ] = 3'd2;
    assign memory3a[85  ] = 3'd2;
    assign memory3a[86  ] = 3'd2;
    assign memory3a[87  ] = 3'd2;
    assign memory3a[88  ] = 3'd0;
    assign memory3a[89  ] = 3'd2;
    assign memory3a[90  ] = 3'd1;
    assign memory3a[91  ] = 3'd2;
    assign memory3a[92  ] = 3'd0;
    assign memory3a[93  ] = 3'd2;
    assign memory3a[94  ] = 3'd2;
    assign memory3a[95  ] = 3'd1;
    assign memory3a[96  ] = 3'd0;
    assign memory3a[97  ] = 3'd2;
    assign memory3a[98  ] = 3'd2;
    assign memory3a[99  ] = 3'd0;
    assign memory3a[100 ] = 3'd2;
    assign memory3a[101 ] = 3'd2;
    assign memory3a[102 ] = 3'd0;
    assign memory3a[103 ] = 3'd1;
    assign memory3a[104 ] = 3'd2;
    assign memory3a[105 ] = 3'd2;
    assign memory3a[106 ] = 3'd2;
    assign memory3a[107 ] = 3'd1;
    assign memory3a[108 ] = 3'd2;
    assign memory3a[109 ] = 3'd2;
    assign memory3a[110 ] = 3'd2;
    assign memory3a[111 ] = 3'd2;
    assign memory3a[112 ] = 3'd2;
    assign memory3a[113 ] = 3'd0;
    assign memory3a[114 ] = 3'd2;
    assign memory3a[115 ] = 3'd1;
    assign memory3a[116 ] = 3'd2;
    assign memory3a[117 ] = 3'd1;
    assign memory3a[118 ] = 3'd2;
    assign memory3a[119 ] = 3'd2;
    assign memory3a[120 ] = 3'd0;
    assign memory3a[121 ] = 3'd2;
    assign memory3a[122 ] = 3'd1;
    assign memory3a[123 ] = 3'd2;
    assign memory3a[124 ] = 3'd0;
    assign memory3a[125 ] = 3'd2;
    assign memory3a[126 ] = 3'd2;
    assign memory3a[127 ] = 3'd1;
    assign memory3a[128 ] = 3'd0;
    assign memory3a[129 ] = 3'd2;
    assign memory3a[130 ] = 3'd0;
    assign memory3a[131 ] = 3'd1;
    assign memory3a[132 ] = 3'd2;
    assign memory3a[133 ] = 3'd2;
    assign memory3a[134 ] = 3'd0;
    assign memory3a[135 ] = 3'd1;
    assign memory3a[136 ] = 3'd2;
    assign memory3a[137 ] = 3'd2;
    assign memory3a[138 ] = 3'd2;
    assign memory3a[139 ] = 3'd1;
    assign memory3a[140 ] = 3'd0;
    assign memory3a[141 ] = 3'd2;
    assign memory3a[142 ] = 3'd2;
    assign memory3a[143 ] = 3'd1;
    assign memory3a[144 ] = 3'd2;
    assign memory3a[145 ] = 3'd0;
    assign memory3a[146 ] = 3'd2;
    assign memory3a[147 ] = 3'd1;
    assign memory3a[148 ] = 3'd2;
    assign memory3a[149 ] = 3'd1;
    assign memory3a[150 ] = 3'd2;
    assign memory3a[151 ] = 3'd2;
    assign memory3a[152 ] = 3'd0;
    assign memory3a[153 ] = 3'd2;
    assign memory3a[154 ] = 3'd1;
    assign memory3a[155 ] = 3'd2;
    assign memory3a[156 ] = 3'd0;
    assign memory3a[157 ] = 3'd2;
    assign memory3a[158 ] = 3'd2;
    assign memory3a[159 ] = 3'd1;
    assign memory3a[160 ] = 3'd0;
    assign memory3a[161 ] = 3'd2;
    assign memory3a[162 ] = 3'd0;
    assign memory3a[163 ] = 3'd1;
    assign memory3a[164 ] = 3'd2;
    assign memory3a[165 ] = 3'd2;
    assign memory3a[166 ] = 3'd0;
    assign memory3a[167 ] = 3'd1;
    assign memory3a[168 ] = 3'd2;
    assign memory3a[169 ] = 3'd2;
    assign memory3a[170 ] = 3'd2;
    assign memory3a[171 ] = 3'd2;
    assign memory3a[172 ] = 3'd0;
    assign memory3a[173 ] = 3'd2;
    assign memory3a[174 ] = 3'd2;
    assign memory3a[175 ] = 3'd1;
    assign memory3a[176 ] = 3'd2;
    assign memory3a[177 ] = 3'd0;
    assign memory3a[178 ] = 3'd2;
    assign memory3a[179 ] = 3'd2;
    assign memory3a[180 ] = 3'd0;
    assign memory3a[181 ] = 3'd1;
    assign memory3a[182 ] = 3'd2;
    assign memory3a[183 ] = 3'd2;
    assign memory3a[184 ] = 3'd0;
    assign memory3a[185 ] = 3'd2;
    assign memory3a[186 ] = 3'd2;
    assign memory3a[187 ] = 3'd2;
    assign memory3a[188 ] = 3'd0;
    assign memory3a[189 ] = 3'd1;
    assign memory3a[190 ] = 3'd2;
    assign memory3a[191 ] = 3'd1;
    assign memory3a[192 ] = 3'd0;
    assign memory3a[193 ] = 3'd2;
    assign memory3a[194 ] = 3'd0;
    assign memory3a[195 ] = 3'd1;
    assign memory3a[196 ] = 3'd0;
    assign memory3a[197 ] = 3'd2;
    assign memory3a[198 ] = 3'd0;
    assign memory3a[199 ] = 3'd1;
    assign memory3a[200 ] = 3'd0;
    assign memory3a[201 ] = 3'd2;
    assign memory3a[202 ] = 3'd2;
    assign memory3a[203 ] = 3'd2;
    assign memory3a[204 ] = 3'd0;
    assign memory3a[205 ] = 3'd2;
    assign memory3a[206 ] = 3'd2;
    assign memory3a[207 ] = 3'd1;
    assign memory3a[208 ] = 3'd2;
    assign memory3a[209 ] = 3'd0;
    assign memory3a[210 ] = 3'd2;
    assign memory3a[211 ] = 3'd2;
    assign memory3a[212 ] = 3'd0;
    assign memory3a[213 ] = 3'd1;
    assign memory3a[214 ] = 3'd2;
    assign memory3a[215 ] = 3'd1;
    assign memory3a[216 ] = 3'd0;
    assign memory3a[217 ] = 3'd2;
    assign memory3a[218 ] = 3'd2;
    assign memory3a[219 ] = 3'd2;
    assign memory3a[220 ] = 3'd0;
    assign memory3a[221 ] = 3'd1;
    assign memory3a[222 ] = 3'd0;
    assign memory3a[223 ] = 3'd2;
    assign memory3a[224 ] = 3'd2;
    assign memory3a[225 ] = 3'd2;
    assign memory3a[226 ] = 3'd0;
    assign memory3a[227 ] = 3'd2;
    assign memory3a[228 ] = 3'd0;
    assign memory3a[229 ] = 3'd2;
    assign memory3a[230 ] = 3'd2;
    assign memory3a[231 ] = 3'd1;
    assign memory3a[232 ] = 3'd0;
    assign memory3a[233 ] = 3'd2;
    assign memory3a[234 ] = 3'd2;
    assign memory3a[235 ] = 3'd2;
    assign memory3a[236 ] = 3'd0;
    assign memory3a[237 ] = 3'd2;
    assign memory3a[238 ] = 3'd0;
    assign memory3a[239 ] = 3'd1;
    assign memory3a[240 ] = 3'd2;
    assign memory3a[241 ] = 3'd2;
    assign memory3a[242 ] = 3'd2;
    assign memory3a[243 ] = 3'd2;
    assign memory3a[244 ] = 3'd0;
    assign memory3a[245 ] = 3'd1;
    assign memory3a[246 ] = 3'd2;
    assign memory3a[247 ] = 3'd1;
    assign memory3a[248 ] = 3'd2;
    assign memory3a[249 ] = 3'd2;
    assign memory3a[250 ] = 3'd2;
    assign memory3a[251 ] = 3'd1;
    assign memory3a[252 ] = 3'd2;
    assign memory3a[253 ] = 3'd1;
    assign memory3a[254 ] = 3'd0;
    assign memory3a[255 ] = 3'd2;
    assign memory3a[256 ] = 3'd2;
    assign memory3a[257 ] = 3'd2;
    assign memory3a[258 ] = 3'd0;
    assign memory3a[259 ] = 3'd2;
    assign memory3a[260 ] = 3'd0;
    assign memory3a[261 ] = 3'd2;
    assign memory3a[262 ] = 3'd2;
    assign memory3a[263 ] = 3'd1;
    assign memory3a[264 ] = 3'd0;
    assign memory3a[265 ] = 3'd1;
    assign memory3a[266 ] = 3'd2;
    assign memory3a[267 ] = 3'd2;
    assign memory3a[268 ] = 3'd0;
    assign memory3a[269 ] = 3'd2;
    assign memory3a[270 ] = 3'd0;
    assign memory3a[271 ] = 3'd1;
    assign memory3a[272 ] = 3'd2;
    assign memory3a[273 ] = 3'd2;
    assign memory3a[274 ] = 3'd2;
    assign memory3a[275 ] = 3'd1;
    assign memory3a[276 ] = 3'd0;
    assign memory3a[277 ] = 3'd2;
    assign memory3a[278 ] = 3'd2;
    assign memory3a[279 ] = 3'd1;
    assign memory3a[280 ] = 3'd2;
    assign memory3a[281 ] = 3'd2;
    assign memory3a[282 ] = 3'd2;
    assign memory3a[283 ] = 3'd1;
    assign memory3a[284 ] = 3'd2;
    assign memory3a[285 ] = 3'd1;
    assign memory3a[286 ] = 3'd0;
    assign memory3a[287 ] = 3'd1;
    assign memory3a[288 ] = 3'd2;
    assign memory3a[289 ] = 3'd1;
    assign memory3a[290 ] = 3'd2;
    assign memory3a[291 ] = 3'd2;
    assign memory3a[292 ] = 3'd0;
    assign memory3a[293 ] = 3'd2;
    assign memory3a[294 ] = 3'd2;
    assign memory3a[295 ] = 3'd2;
    assign memory3a[296 ] = 3'd0;
    assign memory3a[297 ] = 3'd1;
    assign memory3a[298 ] = 3'd2;
    assign memory3a[299 ] = 3'd2;
    assign memory3a[300 ] = 3'd0;
    assign memory3a[301 ] = 3'd2;
    assign memory3a[302 ] = 3'd0;
    assign memory3a[303 ] = 3'd1;
    assign memory3a[304 ] = 3'd2;
    assign memory3a[305 ] = 3'd2;
    assign memory3a[306 ] = 3'd2;
    assign memory3a[307 ] = 3'd1;
    assign memory3a[308 ] = 3'd0;
    assign memory3a[309 ] = 3'd2;
    assign memory3a[310 ] = 3'd2;
    assign memory3a[311 ] = 3'd1;
    assign memory3a[312 ] = 3'd2;
    assign memory3a[313 ] = 3'd3;
    assign memory3a[314 ] = 3'd0;
    assign memory3a[315 ] = 3'd1;
    assign memory3a[316 ] = 3'd2;
    assign memory3a[317 ] = 3'd2;
    assign memory3a[318 ] = 3'd0;
    assign memory3a[319 ] = 3'd1;
    assign memory3a[320 ] = 3'd2;
    assign memory3a[321 ] = 3'd1;
    assign memory3a[322 ] = 3'd2;
    assign memory3a[323 ] = 3'd2;
    assign memory3a[324 ] = 3'd0;
    assign memory3a[325 ] = 3'd2;
    assign memory3a[326 ] = 3'd0;
    assign memory3a[327 ] = 3'd2;
    assign memory3a[328 ] = 3'd2;
    assign memory3a[329 ] = 3'd1;
    assign memory3a[330 ] = 3'd2;
    assign memory3a[331 ] = 3'd0;
    assign memory3a[332 ] = 3'd2;
    assign memory3a[333 ] = 3'd2;
    assign memory3a[334 ] = 3'd0;
    assign memory3a[335 ] = 3'd2;
    assign memory3a[336 ] = 3'd2;
    assign memory3a[337 ] = 3'd2;
    assign memory3a[338 ] = 3'd0;
    assign memory3a[339 ] = 3'd1;
    assign memory3a[340 ] = 3'd2;
    assign memory3a[341 ] = 3'd2;
    assign memory3a[342 ] = 3'd2;
    assign memory3a[343 ] = 3'd1;
    assign memory3a[344 ] = 3'd3;
    assign memory3a[345 ] = 3'd1;
    assign memory3a[346 ] = 3'd0;
    assign memory3a[347 ] = 3'd1;
    assign memory3a[348 ] = 3'd2;
    assign memory3a[349 ] = 3'd2;
    assign memory3a[350 ] = 3'd0;
    assign memory3a[351 ] = 3'd1;
    assign memory3a[352 ] = 3'd2;
    assign memory3a[353 ] = 3'd1;
    assign memory3a[354 ] = 3'd2;
    assign memory3a[355 ] = 3'd2;
    assign memory3a[356 ] = 3'd0;
    assign memory3a[357 ] = 3'd2;
    assign memory3a[358 ] = 3'd0;
    assign memory3a[359 ] = 3'd2;
    assign memory3a[360 ] = 3'd2;
    assign memory3a[361 ] = 3'd1;
    assign memory3a[362 ] = 3'd2;
    assign memory3a[363 ] = 3'd0;
    assign memory3a[364 ] = 3'd2;
    assign memory3a[365 ] = 3'd2;
    assign memory3a[366 ] = 3'd0;
    assign memory3a[367 ] = 3'd2;
    assign memory3a[368 ] = 3'd2;
    assign memory3a[369 ] = 3'd2;
    assign memory3a[370 ] = 3'd3;
    assign memory3a[371 ] = 3'd1;
    assign memory3a[372 ] = 3'd2;
    assign memory3a[373 ] = 3'd2;
    assign memory3a[374 ] = 3'd2;
    assign memory3a[375 ] = 3'd3;
    assign memory3a[376 ] = 3'd2;
    assign memory3a[377 ] = 3'd1;
    assign memory3a[378 ] = 3'd0;
    assign memory3a[379 ] = 3'd1;
    assign memory3a[380 ] = 3'd2;
    assign memory3a[381 ] = 3'd1;
    assign memory3a[382 ] = 3'd0;
    assign memory3a[383 ] = 3'd1;
    assign memory3a[384 ] = 3'd2;
    assign memory3a[385 ] = 3'd1;
    assign memory3a[386 ] = 3'd2;
    assign memory3a[387 ] = 3'd2;
    assign memory3a[388 ] = 3'd0;
    assign memory3a[389 ] = 3'd2;
    assign memory3a[390 ] = 3'd0;
    assign memory3a[391 ] = 3'd2;
    assign memory3a[392 ] = 3'd2;
    assign memory3a[393 ] = 3'd1;
    assign memory3a[394 ] = 3'd2;
    assign memory3a[395 ] = 3'd0;
    assign memory3a[396 ] = 3'd2;
    assign memory3a[397 ] = 3'd2;
    assign memory3a[398 ] = 3'd0;
    assign memory3a[399 ] = 3'd2;
    assign memory3a[400 ] = 3'd2;
    assign memory3a[401 ] = 3'd3;
    assign memory3a[402 ] = 3'd0;
    assign memory3a[403 ] = 3'd1;
    assign memory3a[404 ] = 3'd2;
    assign memory3a[405 ] = 3'd2;
    assign memory3a[406 ] = 3'd2;
    assign memory3a[407 ] = 3'd3;
    assign memory3a[408 ] = 3'd2;
    assign memory3a[409 ] = 3'd1;
    assign memory3a[410 ] = 3'd0;
    assign memory3a[411 ] = 3'd1;
    assign memory3a[412 ] = 3'd2;
    assign memory3a[413 ] = 3'd1;
    assign memory3a[414 ] = 3'd2;
    assign memory3a[415 ] = 3'd1;
    assign memory3a[416 ] = 3'd0;
    assign memory3a[417 ] = 3'd1;
    assign memory3a[418 ] = 3'd2;
    assign memory3a[419 ] = 3'd2;
    assign memory3a[420 ] = 3'd2;
    assign memory3a[421 ] = 3'd2;
    assign memory3a[422 ] = 3'd0;
    assign memory3a[423 ] = 3'd2;
    assign memory3a[424 ] = 3'd2;
    assign memory3a[425 ] = 3'd2;
    assign memory3a[426 ] = 3'd2;
    assign memory3a[427 ] = 3'd0;
    assign memory3a[428 ] = 3'd1;
    assign memory3a[429 ] = 3'd2;
    assign memory3a[430 ] = 3'd0;
    assign memory3a[431 ] = 3'd2;
    assign memory3a[432 ] = 3'd3;
    assign memory3a[433 ] = 3'd2;
    assign memory3a[434 ] = 3'd0;
    assign memory3a[435 ] = 3'd2;
    assign memory3a[436 ] = 3'd2;
    assign memory3a[437 ] = 3'd1;
    assign memory3a[438 ] = 3'd2;
    assign memory3a[439 ] = 3'd3;
    assign memory3a[440 ] = 3'd2;
    assign memory3a[441 ] = 3'd1;
    assign memory3a[442 ] = 3'd0;
    assign memory3a[443 ] = 3'd2;
    assign memory3a[444 ] = 3'd2;
    assign memory3a[445 ] = 3'd1;
    assign memory3a[446 ] = 3'd2;
    assign memory3a[447 ] = 3'd2;
    assign memory3a[448 ] = 3'd0;
    assign memory3a[449 ] = 3'd1;
    assign memory3a[450 ] = 3'd2;
    assign memory3a[451 ] = 3'd2;
    assign memory3a[452 ] = 3'd2;
    assign memory3a[453 ] = 3'd1;
    assign memory3a[454 ] = 3'd0;
    assign memory3a[455 ] = 3'd2;
    assign memory3a[456 ] = 3'd2;
    assign memory3a[457 ] = 3'd2;
    assign memory3a[458 ] = 3'd2;
    assign memory3a[459 ] = 3'd0;
    assign memory3a[460 ] = 3'd1;
    assign memory3a[461 ] = 3'd2;
    assign memory3a[462 ] = 3'd2;
    assign memory3a[463 ] = 3'd2;
    assign memory3a[464 ] = 3'd3;
    assign memory3a[465 ] = 3'd2;
    assign memory3a[466 ] = 3'd0;
    assign memory3a[467 ] = 3'd2;
    assign memory3a[468 ] = 3'd2;
    assign memory3a[469 ] = 3'd1;
    assign memory3a[470 ] = 3'd2;
    assign memory3a[471 ] = 3'd3;
    assign memory3a[472 ] = 3'd2;
    assign memory3a[473 ] = 3'd1;
    assign memory3a[474 ] = 3'd2;
    assign memory3a[475 ] = 3'd2;
    assign memory3a[476 ] = 3'd2;
    assign memory3a[477 ] = 3'd1;
    assign memory3a[478 ] = 3'd2;
    assign memory3a[479 ] = 3'd2;
    assign memory3a[480 ] = 3'd0;
    assign memory3a[481 ] = 3'd2;
    assign memory3a[482 ] = 3'd2;
    assign memory3a[483 ] = 3'd2;
    assign memory3a[484 ] = 3'd2;
    assign memory3a[485 ] = 3'd1;
    assign memory3a[486 ] = 3'd2;
    assign memory3a[487 ] = 3'd2;
    assign memory3a[488 ] = 3'd0;
    assign memory3a[489 ] = 3'd2;
    assign memory3a[490 ] = 3'd2;
    assign memory3a[491 ] = 3'd2;
    assign memory3a[492 ] = 3'd1;
    assign memory3a[493 ] = 3'd2;
    assign memory3a[494 ] = 3'd2;
    assign memory3a[495 ] = 3'd2;
    assign memory3a[496 ] = 3'd3;
    assign memory3a[497 ] = 3'd2;
    assign memory3a[498 ] = 3'd2;
    assign memory3a[499 ] = 3'd2;
    assign memory3a[500 ] = 3'd0;
    assign memory3a[501 ] = 3'd1;
    assign memory3a[502 ] = 3'd2;
    assign memory3a[503 ] = 3'd3;
    assign memory3a[504 ] = 3'd2;
    assign memory3a[505 ] = 3'd2;
    assign memory3a[506 ] = 3'd2;
    assign memory3a[507 ] = 3'd2;
    assign memory3a[508 ] = 3'd2;
    assign memory3a[509 ] = 3'd1;
    assign memory3a[510 ] = 3'd2;
    assign memory3a[511 ] = 3'd2;
    assign memory3a[512 ] = 3'd0;
    assign memory3a[513 ] = 3'd2;
    assign memory3a[514 ] = 3'd2;
    assign memory3a[515 ] = 3'd0;
    assign memory3a[516 ] = 3'd2;
    assign memory3a[517 ] = 3'd1;
    assign memory3a[518 ] = 3'd2;
    assign memory3a[519 ] = 3'd0;
    assign memory3a[520 ] = 3'd2;
    assign memory3a[521 ] = 3'd2;
    assign memory3a[522 ] = 3'd2;
    assign memory3a[523 ] = 3'd2;
    assign memory3a[524 ] = 3'd1;
    assign memory3a[525 ] = 3'd2;
    assign memory3a[526 ] = 3'd2;
    assign memory3a[527 ] = 3'd2;
    assign memory3a[528 ] = 3'd3;
    assign memory3a[529 ] = 3'd1;
    assign memory3a[530 ] = 3'd2;
    assign memory3a[531 ] = 3'd2;
    assign memory3a[532 ] = 3'd0;
    assign memory3a[533 ] = 3'd1;
    assign memory3a[534 ] = 3'd2;
    assign memory3a[535 ] = 3'd2;
    assign memory3a[536 ] = 3'd0;
    assign memory3a[537 ] = 3'd2;
    assign memory3a[538 ] = 3'd2;
    assign memory3a[539 ] = 3'd2;
    assign memory3a[540 ] = 3'd0;
    assign memory3a[541 ] = 3'd1;
    assign memory3a[542 ] = 3'd2;
    assign memory3a[543 ] = 3'd2;
    assign memory3a[544 ] = 3'd0;
    assign memory3a[545 ] = 3'd2;
    assign memory3a[546 ] = 3'd1;
    assign memory3a[547 ] = 3'd0;
    assign memory3a[548 ] = 3'd2;
    assign memory3a[549 ] = 3'd1;
    assign memory3a[550 ] = 3'd2;
    assign memory3a[551 ] = 3'd0;
    assign memory3a[552 ] = 3'd2;
    assign memory3a[553 ] = 3'd0;
    assign memory3a[554 ] = 3'd2;
    assign memory3a[555 ] = 3'd2;
    assign memory3a[556 ] = 3'd1;
    assign memory3a[557 ] = 3'd2;
    assign memory3a[558 ] = 3'd2;
    assign memory3a[559 ] = 3'd2;
    assign memory3a[560 ] = 3'd3;
    assign memory3a[561 ] = 3'd1;
    assign memory3a[562 ] = 3'd2;
    assign memory3a[563 ] = 3'd2;
    assign memory3a[564 ] = 3'd0;
    assign memory3a[565 ] = 3'd1;
    assign memory3a[566 ] = 3'd2;
    assign memory3a[567 ] = 3'd2;
    assign memory3a[568 ] = 3'd0;
    assign memory3a[569 ] = 3'd2;
    assign memory3a[570 ] = 3'd1;
    assign memory3a[571 ] = 3'd2;
    assign memory3a[572 ] = 3'd0;
    assign memory3a[573 ] = 3'd2;
    assign memory3a[574 ] = 3'd2;
    assign memory3a[575 ] = 3'd2;
    assign memory3a[576 ] = 3'd0;
    assign memory3a[577 ] = 3'd2;
    assign memory3a[578 ] = 3'd1;
    assign memory3a[579 ] = 3'd0;
    assign memory3a[580 ] = 3'd2;
    assign memory3a[581 ] = 3'd1;
    assign memory3a[582 ] = 3'd2;
    assign memory3a[583 ] = 3'd0;
    assign memory3a[584 ] = 3'd2;
    assign memory3a[585 ] = 3'd0;
    assign memory3a[586 ] = 3'd2;
    assign memory3a[587 ] = 3'd2;
    assign memory3a[588 ] = 3'd2;
    assign memory3a[589 ] = 3'd2;
    assign memory3a[590 ] = 3'd3;
    assign memory3a[591 ] = 3'd2;
    assign memory3a[592 ] = 3'd3;
    assign memory3a[593 ] = 3'd1;
    assign memory3a[594 ] = 3'd2;
    assign memory3a[595 ] = 3'd2;
    assign memory3a[596 ] = 3'd0;
    assign memory3a[597 ] = 3'd2;
    assign memory3a[598 ] = 3'd2;
    assign memory3a[599 ] = 3'd2;
    assign memory3a[600 ] = 3'd0;
    assign memory3a[601 ] = 3'd2;
    assign memory3a[602 ] = 3'd1;
    assign memory3a[603 ] = 3'd2;
    assign memory3a[604 ] = 3'd0;
    assign memory3a[605 ] = 3'd2;
    assign memory3a[606 ] = 3'd2;
    assign memory3a[607 ] = 3'd2;
    assign memory3a[608 ] = 3'd2;
    assign memory3a[609 ] = 3'd2;
    assign memory3a[610 ] = 3'd1;
    assign memory3a[611 ] = 3'd0;
    assign memory3a[612 ] = 3'd2;
    assign memory3a[613 ] = 3'd1;
    assign memory3a[614 ] = 3'd2;
    assign memory3a[615 ] = 3'd0;
    assign memory3a[616 ] = 3'd2;
    assign memory3a[617 ] = 3'd0;
    assign memory3a[618 ] = 3'd2;
    assign memory3a[619 ] = 3'd2;
    assign memory3a[620 ] = 3'd2;
    assign memory3a[621 ] = 3'd3;
    assign memory3a[622 ] = 3'd2;
    assign memory3a[623 ] = 3'd0;
    assign memory3a[624 ] = 3'd2;
    assign memory3a[625 ] = 3'd1;
    assign memory3a[626 ] = 3'd2;
    assign memory3a[627 ] = 3'd2;
    assign memory3a[628 ] = 3'd0;
    assign memory3a[629 ] = 3'd2;
    assign memory3a[630 ] = 3'd2;
    assign memory3a[631 ] = 3'd2;
    assign memory3a[632 ] = 3'd0;
    assign memory3a[633 ] = 3'd2;
    assign memory3a[634 ] = 3'd1;
    assign memory3a[635 ] = 3'd2;
    assign memory3a[636 ] = 3'd0;
    assign memory3a[637 ] = 3'd1;
    assign memory3a[638 ] = 3'd2;
    assign memory3a[639 ] = 3'd2;
    assign memory3a[640 ] = 3'd2;
    assign memory3a[641 ] = 3'd2;
    assign memory3a[642 ] = 3'd1;
    assign memory3a[643 ] = 3'd0;
    assign memory3a[644 ] = 3'd2;
    assign memory3a[645 ] = 3'd2;
    assign memory3a[646 ] = 3'd2;
    assign memory3a[647 ] = 3'd0;
    assign memory3a[648 ] = 3'd2;
    assign memory3a[649 ] = 3'd0;
    assign memory3a[650 ] = 3'd1;
    assign memory3a[651 ] = 3'd0;
    assign memory3a[652 ] = 3'd3;
    assign memory3a[653 ] = 3'd2;
    assign memory3a[654 ] = 3'd2;
    assign memory3a[655 ] = 3'd0;
    assign memory3a[656 ] = 3'd2;
    assign memory3a[657 ] = 3'd1;
    assign memory3a[658 ] = 3'd2;
    assign memory3a[659 ] = 3'd2;
    assign memory3a[660 ] = 3'd2;
    assign memory3a[661 ] = 3'd2;
    assign memory3a[662 ] = 3'd2;
    assign memory3a[663 ] = 3'd1;
    assign memory3a[664 ] = 3'd0;
    assign memory3a[665 ] = 3'd2;
    assign memory3a[666 ] = 3'd1;
    assign memory3a[667 ] = 3'd2;
    assign memory3a[668 ] = 3'd0;
    assign memory3a[669 ] = 3'd1;
    assign memory3a[670 ] = 3'd2;
    assign memory3a[671 ] = 3'd2;
    assign memory3a[672 ] = 3'd2;
    assign memory3a[673 ] = 3'd0;
    assign memory3a[674 ] = 3'd1;
    assign memory3a[675 ] = 3'd0;
    assign memory3a[676 ] = 3'd2;
    assign memory3a[677 ] = 3'd2;
    assign memory3a[678 ] = 3'd2;
    assign memory3a[679 ] = 3'd0;
    assign memory3a[680 ] = 3'd2;
    assign memory3a[681 ] = 3'd0;
    assign memory3a[682 ] = 3'd1;
    assign memory3a[683 ] = 3'd0;
    assign memory3a[684 ] = 3'd3;
    assign memory3a[685 ] = 3'd2;
    assign memory3a[686 ] = 3'd1;
    assign memory3a[687 ] = 3'd0;
    assign memory3a[688 ] = 3'd2;
    assign memory3a[689 ] = 3'd1;
    assign memory3a[690 ] = 3'd2;
    assign memory3a[691 ] = 3'd2;
    assign memory3a[692 ] = 3'd1;
    assign memory3a[693 ] = 3'd2;
    assign memory3a[694 ] = 3'd0;
    assign memory3a[695 ] = 3'd1;
    assign memory3a[696 ] = 3'd2;
    assign memory3a[697 ] = 3'd2;
    assign memory3a[698 ] = 3'd1;
    assign memory3a[699 ] = 3'd2;
    assign memory3a[700 ] = 3'd2;
    assign memory3a[701 ] = 3'd1;
    assign memory3a[702 ] = 3'd2;
    assign memory3a[703 ] = 3'd1;
    assign memory3a[704 ] = 3'd2;
    assign memory3a[705 ] = 3'd0;
    assign memory3a[706 ] = 3'd2;
    assign memory3a[707 ] = 3'd2;
    assign memory3a[708 ] = 3'd2;
    assign memory3a[709 ] = 3'd2;
    assign memory3a[710 ] = 3'd2;
    assign memory3a[711 ] = 3'd2;
    assign memory3a[712 ] = 3'd2;
    assign memory3a[713 ] = 3'd2;
    assign memory3a[714 ] = 3'd1;
    assign memory3a[715 ] = 3'd0;
    assign memory3a[716 ] = 3'd3;
    assign memory3a[717 ] = 3'd2;
    assign memory3a[718 ] = 3'd1;
    assign memory3a[719 ] = 3'd0;
    assign memory3a[720 ] = 3'd2;
    assign memory3a[721 ] = 3'd1;
    assign memory3a[722 ] = 3'd0;
    assign memory3a[723 ] = 3'd2;
    assign memory3a[724 ] = 3'd1;
    assign memory3a[725 ] = 3'd2;
    assign memory3a[726 ] = 3'd0;
    assign memory3a[727 ] = 3'd1;
    assign memory3a[728 ] = 3'd2;
    assign memory3a[729 ] = 3'd2;
    assign memory3a[730 ] = 3'd2;
    assign memory3a[731 ] = 3'd2;
    assign memory3a[732 ] = 3'd2;
    assign memory3a[733 ] = 3'd1;
    assign memory3a[734 ] = 3'd2;
    assign memory3a[735 ] = 3'd1;
    assign memory3a[736 ] = 3'd2;
    assign memory3a[737 ] = 3'd0;
    assign memory3a[738 ] = 3'd2;
    assign memory3a[739 ] = 3'd2;
    assign memory3a[740 ] = 3'd2;
    assign memory3a[741 ] = 3'd2;
    assign memory3a[742 ] = 3'd0;
    assign memory3a[743 ] = 3'd2;
    assign memory3a[744 ] = 3'd2;
    assign memory3a[745 ] = 3'd2;
    assign memory3a[746 ] = 3'd1;
    assign memory3a[747 ] = 3'd0;
    assign memory3a[748 ] = 3'd3;
    assign memory3a[749 ] = 3'd2;
    assign memory3a[750 ] = 3'd1;
    assign memory3a[751 ] = 3'd0;
    assign memory3a[752 ] = 3'd2;
    assign memory3a[753 ] = 3'd2;
    assign memory3a[754 ] = 3'd0;
    assign memory3a[755 ] = 3'd2;
    assign memory3a[756 ] = 3'd1;
    assign memory3a[757 ] = 3'd2;
    assign memory3a[758 ] = 3'd0;
    assign memory3a[759 ] = 3'd1;
    assign memory3a[760 ] = 3'd2;
    assign memory3a[761 ] = 3'd2;
    assign memory3a[762 ] = 3'd2;
    assign memory3a[763 ] = 3'd2;
    assign memory3a[764 ] = 3'd2;
    assign memory3a[765 ] = 3'd1;
    assign memory3a[766 ] = 3'd2;
    assign memory3a[767 ] = 3'd1;
    assign memory3a[768 ] = 3'd2;
    assign memory3a[769 ] = 3'd0;
    assign memory3a[770 ] = 3'd2;
    assign memory3a[771 ] = 3'd2;
    assign memory3a[772 ] = 3'd2;
    assign memory3a[773 ] = 3'd0;
    assign memory3a[774 ] = 3'd2;
    assign memory3a[775 ] = 3'd1;
    assign memory3a[776 ] = 3'd2;
    assign memory3a[777 ] = 3'd2;
    assign memory3a[778 ] = 3'd1;
    assign memory3a[779 ] = 3'd0;
    assign memory3a[780 ] = 3'd3;
    assign memory3a[781 ] = 3'd2;
    assign memory3a[782 ] = 3'd1;
    assign memory3a[783 ] = 3'd0;
    assign memory3a[784 ] = 3'd2;
    assign memory3a[785 ] = 3'd2;
    assign memory3a[786 ] = 3'd0;
    assign memory3a[787 ] = 3'd2;
    assign memory3a[788 ] = 3'd1;
    assign memory3a[789 ] = 3'd2;
    assign memory3a[790 ] = 3'd0;
    assign memory3a[791 ] = 3'd1;
    assign memory3a[792 ] = 3'd2;
    assign memory3a[793 ] = 3'd2;
    assign memory3a[794 ] = 3'd3;
    assign memory3a[795 ] = 3'd1;
    assign memory3a[796 ] = 3'd2;
    assign memory3a[797 ] = 3'd2;
    assign memory3a[798 ] = 3'd2;
    assign memory3a[799 ] = 3'd1;
    assign memory3a[800 ] = 3'd2;
    assign memory3a[801 ] = 3'd0;
    assign memory3a[802 ] = 3'd2;
    assign memory3a[803 ] = 3'd2;
    assign memory3a[804 ] = 3'd2;
    assign memory3a[805 ] = 3'd0;
    assign memory3a[806 ] = 3'd2;
    assign memory3a[807 ] = 3'd1;
    assign memory3a[808 ] = 3'd2;
    assign memory3a[809 ] = 3'd0;
    assign memory3a[810 ] = 3'd1;
    assign memory3a[811 ] = 3'd2;
    assign memory3a[812 ] = 3'd3;
    assign memory3a[813 ] = 3'd2;
    assign memory3a[814 ] = 3'd1;
    assign memory3a[815 ] = 3'd2;
    assign memory3a[816 ] = 3'd2;
    assign memory3a[817 ] = 3'd2;
    assign memory3a[818 ] = 3'd0;
    assign memory3a[819 ] = 3'd2;
    assign memory3a[820 ] = 3'd1;
    assign memory3a[821 ] = 3'd2;
    assign memory3a[822 ] = 3'd0;
    assign memory3a[823 ] = 3'd1;
    assign memory3a[824 ] = 3'd2;
    assign memory3a[825 ] = 3'd3;
    assign memory3a[826 ] = 3'd0;
    assign memory3a[827 ] = 3'd1;
    assign memory3a[828 ] = 3'd2;
    assign memory3a[829 ] = 3'd2;
    assign memory3a[830 ] = 3'd2;
    assign memory3a[831 ] = 3'd1;
    assign memory3a[832 ] = 3'd2;
    assign memory3a[833 ] = 3'd2;
    assign memory3a[834 ] = 3'd2;
    assign memory3a[835 ] = 3'd0;
    assign memory3a[836 ] = 3'd2;
    assign memory3a[837 ] = 3'd0;
    assign memory3a[838 ] = 3'd2;
    assign memory3a[839 ] = 3'd1;
    assign memory3a[840 ] = 3'd0;
    assign memory3a[841 ] = 3'd2;
    assign memory3a[842 ] = 3'd2;
    assign memory3a[843 ] = 3'd2;
    assign memory3a[844 ] = 3'd2;
    assign memory3a[845 ] = 3'd0;
    assign memory3a[846 ] = 3'd2;
    assign memory3a[847 ] = 3'd2;
    assign memory3a[848 ] = 3'd2;
    assign memory3a[849 ] = 3'd2;
    assign memory3a[850 ] = 3'd2;
    assign memory3a[851 ] = 3'd2;
    assign memory3a[852 ] = 3'd1;
    assign memory3a[853 ] = 3'd2;
    assign memory3a[854 ] = 3'd2;
    assign memory3a[855 ] = 3'd2;
    assign memory3a[856 ] = 3'd3;
    assign memory3a[857 ] = 3'd2;
    assign memory3a[858 ] = 3'd0;
    assign memory3a[859 ] = 3'd1;
    assign memory3a[860 ] = 3'd2;
    assign memory3a[861 ] = 3'd2;
    assign memory3a[862 ] = 3'd2;
    assign memory3a[863 ] = 3'd1;
    assign memory3a[864 ] = 3'd2;
    assign memory3a[865 ] = 3'd2;
    assign memory3a[866 ] = 3'd0;
    assign memory3a[867 ] = 3'd2;
    assign memory3a[868 ] = 3'd2;
    assign memory3a[869 ] = 3'd0;
    assign memory3a[870 ] = 3'd2;
    assign memory3a[871 ] = 3'd1;
    assign memory3a[872 ] = 3'd0;
    assign memory3a[873 ] = 3'd2;
    assign memory3a[874 ] = 3'd2;
    assign memory3a[875 ] = 3'd2;
    assign memory3a[876 ] = 3'd0;
    assign memory3a[877 ] = 3'd2;
    assign memory3a[878 ] = 3'd2;
    assign memory3a[879 ] = 3'd2;
    assign memory3a[880 ] = 3'd2;
    assign memory3a[881 ] = 3'd2;
    assign memory3a[882 ] = 3'd2;
    assign memory3a[883 ] = 3'd2;
    assign memory3a[884 ] = 3'd2;
    assign memory3a[885 ] = 3'd2;
    assign memory3a[886 ] = 3'd2;
    assign memory3a[887 ] = 3'd0;
    assign memory3a[888 ] = 3'd3;
    assign memory3a[889 ] = 3'd2;
    assign memory3a[890 ] = 3'd0;
    assign memory3a[891 ] = 3'd1;
    assign memory3a[892 ] = 3'd2;
    assign memory3a[893 ] = 3'd2;
    assign memory3a[894 ] = 3'd2;
    assign memory3a[895 ] = 3'd2;
    assign memory3a[896 ] = 3'd2;
    assign memory3a[897 ] = 3'd2;
    assign memory3a[898 ] = 3'd0;
    assign memory3a[899 ] = 3'd2;
    assign memory3a[900 ] = 3'd1;
    assign memory3a[901 ] = 3'd0;
    assign memory3a[902 ] = 3'd2;
    assign memory3a[903 ] = 3'd1;
    assign memory3a[904 ] = 3'd0;
    assign memory3a[905 ] = 3'd2;
    assign memory3a[906 ] = 3'd2;
    assign memory3a[907 ] = 3'd2;
    assign memory3a[908 ] = 3'd0;
    assign memory3a[909 ] = 3'd2;
    assign memory3a[910 ] = 3'd2;
    assign memory3a[911 ] = 3'd1;
    assign memory3a[912 ] = 3'd2;
    assign memory3a[913 ] = 3'd2;
    assign memory3a[914 ] = 3'd1;
    assign memory3a[915 ] = 3'd2;
    assign memory3a[916 ] = 3'd2;
    assign memory3a[917 ] = 3'd2;
    assign memory3a[918 ] = 3'd0;
    assign memory3a[919 ] = 3'd2;
    assign memory3a[920 ] = 3'd3;
    assign memory3a[921 ] = 3'd1;
    assign memory3a[922 ] = 3'd0;
    assign memory3a[923 ] = 3'd1;
    assign memory3a[924 ] = 3'd2;
    assign memory3a[925 ] = 3'd2;
    assign memory3a[926 ] = 3'd2;
    assign memory3a[927 ] = 3'd2;
    assign memory3a[928 ] = 3'd0;
    assign memory3a[929 ] = 3'd2;
    assign memory3a[930 ] = 3'd0;
    assign memory3a[931 ] = 3'd2;
    assign memory3a[932 ] = 3'd1;
    assign memory3a[933 ] = 3'd2;
    assign memory3a[934 ] = 3'd2;
    assign memory3a[935 ] = 3'd1;
    assign memory3a[936 ] = 3'd0;
    assign memory3a[937 ] = 3'd2;
    assign memory3a[938 ] = 3'd0;
    assign memory3a[939 ] = 3'd2;
    assign memory3a[940 ] = 3'd0;
    assign memory3a[941 ] = 3'd2;
    assign memory3a[942 ] = 3'd1;
    assign memory3a[943 ] = 3'd2;
    assign memory3a[944 ] = 3'd2;
    assign memory3a[945 ] = 3'd2;
    assign memory3a[946 ] = 3'd1;
    assign memory3a[947 ] = 3'd2;
    assign memory3a[948 ] = 3'd2;
    assign memory3a[949 ] = 3'd0;
    assign memory3a[950 ] = 3'd2;
    assign memory3a[951 ] = 3'd2;
    assign memory3a[952 ] = 3'd3;
    assign memory3a[953 ] = 3'd1;
    assign memory3a[954 ] = 3'd0;
    assign memory3a[955 ] = 3'd2;
    assign memory3a[956 ] = 3'd2;
    assign memory3a[957 ] = 3'd2;
    assign memory3a[958 ] = 3'd2;
    assign memory3a[959 ] = 3'd2;
    assign memory3a[960 ] = 3'd0;
    assign memory3a[961 ] = 3'd2;
    assign memory3a[962 ] = 3'd0;
    assign memory3a[963 ] = 3'd2;
    assign memory3a[964 ] = 3'd1;
    assign memory3a[965 ] = 3'd2;
    assign memory3a[966 ] = 3'd2;
    assign memory3a[967 ] = 3'd1;
    assign memory3a[968 ] = 3'd0;
    assign memory3a[969 ] = 3'd2;
    assign memory3a[970 ] = 3'd0;
    assign memory3a[971 ] = 3'd2;
    assign memory3a[972 ] = 3'd0;
    assign memory3a[973 ] = 3'd1;
    assign memory3a[974 ] = 3'd2;
    assign memory3a[975 ] = 3'd2;
    assign memory3a[976 ] = 3'd2;
    assign memory3a[977 ] = 3'd2;
    assign memory3a[978 ] = 3'd1;
    assign memory3a[979 ] = 3'd2;
    assign memory3a[980 ] = 3'd2;
    assign memory3a[981 ] = 3'd0;
    assign memory3a[982 ] = 3'd2;
    assign memory3a[983 ] = 3'd2;
    assign memory3a[984 ] = 3'd3;
    assign memory3a[985 ] = 3'd1;
    assign memory3a[986 ] = 3'd2;
    assign memory3a[987 ] = 3'd2;
    assign memory3a[988 ] = 3'd2;
    assign memory3a[989 ] = 3'd2;
    assign memory3a[990 ] = 3'd2;
    assign memory3a[991 ] = 3'd2;
    assign memory3a[992 ] = 3'd0;
    assign memory3a[993 ] = 3'd2;
    assign memory3a[994 ] = 3'd0;
    assign memory3a[995 ] = 3'd2;
    assign memory3a[996 ] = 3'd1;
    assign memory3a[997 ] = 3'd2;
    assign memory3a[998 ] = 3'd2;
    assign memory3a[999 ] = 3'd2;
    assign memory3a[1000] = 3'd0;
    assign memory3a[1001] = 3'd2;
    assign memory3a[1002] = 3'd0;
    assign memory3a[1003] = 3'd2;
    assign memory3a[1004] = 3'd0;
    assign memory3a[1005] = 3'd1;
    assign memory3a[1006] = 3'd2;
    assign memory3a[1007] = 3'd2;
    assign memory3a[1008] = 3'd2;
    assign memory3a[1009] = 3'd2;
    assign memory3a[1010] = 3'd1;
    assign memory3a[1011] = 3'd2;
    assign memory3a[1012] = 3'd2;
    assign memory3a[1013] = 3'd0;
    assign memory3a[1014] = 3'd2;
    assign memory3a[1015] = 3'd2;
    assign memory3a[1016] = 3'd2;
    assign memory3a[1017] = 3'd1;
    assign memory3a[1018] = 3'd2;
    assign memory3a[1019] = 3'd2;
    assign memory3a[1020] = 3'd2;
    assign memory3a[1021] = 3'd2;
    assign memory3a[1022] = 3'd2;
    assign memory3a[1023] = 3'd2;

    assign memory3b[0   ] = 3'd0;
    assign memory3b[1   ] = 3'd0;
    assign memory3b[2   ] = 3'd0;
    assign memory3b[3   ] = 3'd0;
    assign memory3b[4   ] = 3'd0;
    assign memory3b[5   ] = 3'd0;
    assign memory3b[6   ] = 3'd0;
    assign memory3b[7   ] = 3'd0;
    assign memory3b[8   ] = 3'd0;
    assign memory3b[9   ] = 3'd0;
    assign memory3b[10  ] = 3'd0;
    assign memory3b[11  ] = 3'd0;
    assign memory3b[12  ] = 3'd1;
    assign memory3b[13  ] = 3'd2;
    assign memory3b[14  ] = 3'd0;
    assign memory3b[15  ] = 3'd0;
    assign memory3b[16  ] = 3'd0;
    assign memory3b[17  ] = 3'd0;
    assign memory3b[18  ] = 3'd0;
    assign memory3b[19  ] = 3'd1;
    assign memory3b[20  ] = 3'd0;
    assign memory3b[21  ] = 3'd0;
    assign memory3b[22  ] = 3'd0;
    assign memory3b[23  ] = 3'd0;
    assign memory3b[24  ] = 3'd0;
    assign memory3b[25  ] = 3'd0;
    assign memory3b[26  ] = 3'd0;
    assign memory3b[27  ] = 3'd0;
    assign memory3b[28  ] = 3'd0;
    assign memory3b[29  ] = 3'd0;
    assign memory3b[30  ] = 3'd0;
    assign memory3b[31  ] = 3'd0;
    assign memory3b[32  ] = 3'd0;
    assign memory3b[33  ] = 3'd0;
    assign memory3b[34  ] = 3'd1;
    assign memory3b[35  ] = 3'd0;
    assign memory3b[36  ] = 3'd3;
    assign memory3b[37  ] = 3'd0;
    assign memory3b[38  ] = 3'd0;
    assign memory3b[39  ] = 3'd1;
    assign memory3b[40  ] = 3'd2;
    assign memory3b[41  ] = 3'd3;
    assign memory3b[42  ] = 3'd0;
    assign memory3b[43  ] = 3'd0;
    assign memory3b[44  ] = 3'd0;
    assign memory3b[45  ] = 3'd2;
    assign memory3b[46  ] = 3'd1;
    assign memory3b[47  ] = 3'd0;
    assign memory3b[48  ] = 3'd0;
    assign memory3b[49  ] = 3'd0;
    assign memory3b[50  ] = 3'd3;
    assign memory3b[51  ] = 3'd0;
    assign memory3b[52  ] = 3'd0;
    assign memory3b[53  ] = 3'd3;
    assign memory3b[54  ] = 3'd0;
    assign memory3b[55  ] = 3'd3;
    assign memory3b[56  ] = 3'd0;
    assign memory3b[57  ] = 3'd3;
    assign memory3b[58  ] = 3'd0;
    assign memory3b[59  ] = 3'd0;
    assign memory3b[60  ] = 3'd1;
    assign memory3b[61  ] = 3'd0;
    assign memory3b[62  ] = 3'd0;
    assign memory3b[63  ] = 3'd0;
    assign memory3b[64  ] = 3'd0;
    assign memory3b[65  ] = 3'd0;
    assign memory3b[66  ] = 3'd0;
    assign memory3b[67  ] = 3'd1;
    assign memory3b[68  ] = 3'd0;
    assign memory3b[69  ] = 3'd0;
    assign memory3b[70  ] = 3'd0;
    assign memory3b[71  ] = 3'd0;
    assign memory3b[72  ] = 3'd0;
    assign memory3b[73  ] = 3'd0;
    assign memory3b[74  ] = 3'd0;
    assign memory3b[75  ] = 3'd0;
    assign memory3b[76  ] = 3'd0;
    assign memory3b[77  ] = 3'd0;
    assign memory3b[78  ] = 3'd0;
    assign memory3b[79  ] = 3'd3;
    assign memory3b[80  ] = 3'd0;
    assign memory3b[81  ] = 3'd0;
    assign memory3b[82  ] = 3'd1;
    assign memory3b[83  ] = 3'd1;
    assign memory3b[84  ] = 3'd0;
    assign memory3b[85  ] = 3'd0;
    assign memory3b[86  ] = 3'd2;
    assign memory3b[87  ] = 3'd0;
    assign memory3b[88  ] = 3'd3;
    assign memory3b[89  ] = 3'd0;
    assign memory3b[90  ] = 3'd0;
    assign memory3b[91  ] = 3'd0;
    assign memory3b[92  ] = 3'd0;
    assign memory3b[93  ] = 3'd0;
    assign memory3b[94  ] = 3'd0;
    assign memory3b[95  ] = 3'd0;
    assign memory3b[96  ] = 3'd0;
    assign memory3b[97  ] = 3'd0;
    assign memory3b[98  ] = 3'd3;
    assign memory3b[99  ] = 3'd3;
    assign memory3b[100 ] = 3'd1;
    assign memory3b[101 ] = 3'd0;
    assign memory3b[102 ] = 3'd0;
    assign memory3b[103 ] = 3'd0;
    assign memory3b[104 ] = 3'd0;
    assign memory3b[105 ] = 3'd0;
    assign memory3b[106 ] = 3'd0;
    assign memory3b[107 ] = 3'd0;
    assign memory3b[108 ] = 3'd3;
    assign memory3b[109 ] = 3'd0;
    assign memory3b[110 ] = 3'd0;
    assign memory3b[111 ] = 3'd1;
    assign memory3b[112 ] = 3'd0;
    assign memory3b[113 ] = 3'd3;
    assign memory3b[114 ] = 3'd2;
    assign memory3b[115 ] = 3'd1;
    assign memory3b[116 ] = 3'd0;
    assign memory3b[117 ] = 3'd0;
    assign memory3b[118 ] = 3'd0;
    assign memory3b[119 ] = 3'd0;
    assign memory3b[120 ] = 3'd0;
    assign memory3b[121 ] = 3'd0;
    assign memory3b[122 ] = 3'd0;
    assign memory3b[123 ] = 3'd0;
    assign memory3b[124 ] = 3'd0;
    assign memory3b[125 ] = 3'd0;
    assign memory3b[126 ] = 3'd2;
    assign memory3b[127 ] = 3'd0;
    assign memory3b[128 ] = 3'd0;
    assign memory3b[129 ] = 3'd0;
    assign memory3b[130 ] = 3'd0;
    assign memory3b[131 ] = 3'd3;
    assign memory3b[132 ] = 3'd0;
    assign memory3b[133 ] = 3'd3;
    assign memory3b[134 ] = 3'd0;
    assign memory3b[135 ] = 3'd0;
    assign memory3b[136 ] = 3'd0;
    assign memory3b[137 ] = 3'd0;
    assign memory3b[138 ] = 3'd0;
    assign memory3b[139 ] = 3'd0;
    assign memory3b[140 ] = 3'd0;
    assign memory3b[141 ] = 3'd0;
    assign memory3b[142 ] = 3'd0;
    assign memory3b[143 ] = 3'd0;
    assign memory3b[144 ] = 3'd0;
    assign memory3b[145 ] = 3'd0;
    assign memory3b[146 ] = 3'd0;
    assign memory3b[147 ] = 3'd0;
    assign memory3b[148 ] = 3'd0;
    assign memory3b[149 ] = 3'd0;
    assign memory3b[150 ] = 3'd3;
    assign memory3b[151 ] = 3'd1;
    assign memory3b[152 ] = 3'd0;
    assign memory3b[153 ] = 3'd0;
    assign memory3b[154 ] = 3'd0;
    assign memory3b[155 ] = 3'd0;
    assign memory3b[156 ] = 3'd0;
    assign memory3b[157 ] = 3'd0;
    assign memory3b[158 ] = 3'd0;
    assign memory3b[159 ] = 3'd0;
    assign memory3b[160 ] = 3'd0;
    assign memory3b[161 ] = 3'd3;
    assign memory3b[162 ] = 3'd0;
    assign memory3b[163 ] = 3'd3;
    assign memory3b[164 ] = 3'd0;
    assign memory3b[165 ] = 3'd0;
    assign memory3b[166 ] = 3'd0;
    assign memory3b[167 ] = 3'd0;
    assign memory3b[168 ] = 3'd0;
    assign memory3b[169 ] = 3'd0;
    assign memory3b[170 ] = 3'd3;
    assign memory3b[171 ] = 3'd0;
    assign memory3b[172 ] = 3'd0;
    assign memory3b[173 ] = 3'd0;
    assign memory3b[174 ] = 3'd0;
    assign memory3b[175 ] = 3'd0;
    assign memory3b[176 ] = 3'd3;
    assign memory3b[177 ] = 3'd0;
    assign memory3b[178 ] = 3'd1;
    assign memory3b[179 ] = 3'd0;
    assign memory3b[180 ] = 3'd0;
    assign memory3b[181 ] = 3'd3;
    assign memory3b[182 ] = 3'd0;
    assign memory3b[183 ] = 3'd1;
    assign memory3b[184 ] = 3'd0;
    assign memory3b[185 ] = 3'd0;
    assign memory3b[186 ] = 3'd0;
    assign memory3b[187 ] = 3'd0;
    assign memory3b[188 ] = 3'd0;
    assign memory3b[189 ] = 3'd0;
    assign memory3b[190 ] = 3'd0;
    assign memory3b[191 ] = 3'd0;
    assign memory3b[192 ] = 3'd0;
    assign memory3b[193 ] = 3'd0;
    assign memory3b[194 ] = 3'd0;
    assign memory3b[195 ] = 3'd0;
    assign memory3b[196 ] = 3'd1;
    assign memory3b[197 ] = 3'd0;
    assign memory3b[198 ] = 3'd0;
    assign memory3b[199 ] = 3'd0;
    assign memory3b[200 ] = 3'd0;
    assign memory3b[201 ] = 3'd0;
    assign memory3b[202 ] = 3'd0;
    assign memory3b[203 ] = 3'd0;
    assign memory3b[204 ] = 3'd2;
    assign memory3b[205 ] = 3'd1;
    assign memory3b[206 ] = 3'd0;
    assign memory3b[207 ] = 3'd0;
    assign memory3b[208 ] = 3'd0;
    assign memory3b[209 ] = 3'd0;
    assign memory3b[210 ] = 3'd0;
    assign memory3b[211 ] = 3'd3;
    assign memory3b[212 ] = 3'd0;
    assign memory3b[213 ] = 3'd4;
    assign memory3b[214 ] = 3'd5;
    assign memory3b[215 ] = 3'd0;
    assign memory3b[216 ] = 3'd0;
    assign memory3b[217 ] = 3'd0;
    assign memory3b[218 ] = 3'd0;
    assign memory3b[219 ] = 3'd1;
    assign memory3b[220 ] = 3'd0;
    assign memory3b[221 ] = 3'd0;
    assign memory3b[222 ] = 3'd0;
    assign memory3b[223 ] = 3'd0;
    assign memory3b[224 ] = 3'd0;
    assign memory3b[225 ] = 3'd0;
    assign memory3b[226 ] = 3'd0;
    assign memory3b[227 ] = 3'd0;
    assign memory3b[228 ] = 3'd3;
    assign memory3b[229 ] = 3'd0;
    assign memory3b[230 ] = 3'd0;
    assign memory3b[231 ] = 3'd0;
    assign memory3b[232 ] = 3'd0;
    assign memory3b[233 ] = 3'd2;
    assign memory3b[234 ] = 3'd0;
    assign memory3b[235 ] = 3'd3;
    assign memory3b[236 ] = 3'd1;
    assign memory3b[237 ] = 3'd0;
    assign memory3b[238 ] = 3'd0;
    assign memory3b[239 ] = 3'd0;
    assign memory3b[240 ] = 3'd3;
    assign memory3b[241 ] = 3'd0;
    assign memory3b[242 ] = 3'd1;
    assign memory3b[243 ] = 3'd0;
    assign memory3b[244 ] = 3'd4;
    assign memory3b[245 ] = 3'd4;
    assign memory3b[246 ] = 3'd4;
    assign memory3b[247 ] = 3'd5;
    assign memory3b[248 ] = 3'd3;
    assign memory3b[249 ] = 3'd0;
    assign memory3b[250 ] = 3'd0;
    assign memory3b[251 ] = 3'd0;
    assign memory3b[252 ] = 3'd0;
    assign memory3b[253 ] = 3'd0;
    assign memory3b[254 ] = 3'd0;
    assign memory3b[255 ] = 3'd0;
    assign memory3b[256 ] = 3'd0;
    assign memory3b[257 ] = 3'd0;
    assign memory3b[258 ] = 3'd0;
    assign memory3b[259 ] = 3'd2;
    assign memory3b[260 ] = 3'd0;
    assign memory3b[261 ] = 3'd0;
    assign memory3b[262 ] = 3'd0;
    assign memory3b[263 ] = 3'd0;
    assign memory3b[264 ] = 3'd0;
    assign memory3b[265 ] = 3'd0;
    assign memory3b[266 ] = 3'd2;
    assign memory3b[267 ] = 3'd1;
    assign memory3b[268 ] = 3'd0;
    assign memory3b[269 ] = 3'd0;
    assign memory3b[270 ] = 3'd0;
    assign memory3b[271 ] = 3'd3;
    assign memory3b[272 ] = 3'd3;
    assign memory3b[273 ] = 3'd0;
    assign memory3b[274 ] = 3'd0;
    assign memory3b[275 ] = 3'd0;
    assign memory3b[276 ] = 3'd4;
    assign memory3b[277 ] = 3'd4;
    assign memory3b[278 ] = 3'd4;
    assign memory3b[279 ] = 3'd5;
    assign memory3b[280 ] = 3'd5;
    assign memory3b[281 ] = 3'd3;
    assign memory3b[282 ] = 3'd0;
    assign memory3b[283 ] = 3'd0;
    assign memory3b[284 ] = 3'd0;
    assign memory3b[285 ] = 3'd0;
    assign memory3b[286 ] = 3'd0;
    assign memory3b[287 ] = 3'd0;
    assign memory3b[288 ] = 3'd0;
    assign memory3b[289 ] = 3'd3;
    assign memory3b[290 ] = 3'd0;
    assign memory3b[291 ] = 3'd1;
    assign memory3b[292 ] = 3'd0;
    assign memory3b[293 ] = 3'd0;
    assign memory3b[294 ] = 3'd0;
    assign memory3b[295 ] = 3'd0;
    assign memory3b[296 ] = 3'd0;
    assign memory3b[297 ] = 3'd0;
    assign memory3b[298 ] = 3'd0;
    assign memory3b[299 ] = 3'd1;
    assign memory3b[300 ] = 3'd0;
    assign memory3b[301 ] = 3'd2;
    assign memory3b[302 ] = 3'd0;
    assign memory3b[303 ] = 3'd0;
    assign memory3b[304 ] = 3'd6;
    assign memory3b[305 ] = 3'd0;
    assign memory3b[306 ] = 3'd0;
    assign memory3b[307 ] = 3'd4;
    assign memory3b[308 ] = 3'd4;
    assign memory3b[309 ] = 3'd4;
    assign memory3b[310 ] = 3'd4;
    assign memory3b[311 ] = 3'd5;
    assign memory3b[312 ] = 3'd5;
    assign memory3b[313 ] = 3'd0;
    assign memory3b[314 ] = 3'd0;
    assign memory3b[315 ] = 3'd0;
    assign memory3b[316 ] = 3'd1;
    assign memory3b[317 ] = 3'd0;
    assign memory3b[318 ] = 3'd0;
    assign memory3b[319 ] = 3'd1;
    assign memory3b[320 ] = 3'd0;
    assign memory3b[321 ] = 3'd0;
    assign memory3b[322 ] = 3'd0;
    assign memory3b[323 ] = 3'd0;
    assign memory3b[324 ] = 3'd0;
    assign memory3b[325 ] = 3'd0;
    assign memory3b[326 ] = 3'd0;
    assign memory3b[327 ] = 3'd0;
    assign memory3b[328 ] = 3'd0;
    assign memory3b[329 ] = 3'd0;
    assign memory3b[330 ] = 3'd0;
    assign memory3b[331 ] = 3'd3;
    assign memory3b[332 ] = 3'd0;
    assign memory3b[333 ] = 3'd0;
    assign memory3b[334 ] = 3'd0;
    assign memory3b[335 ] = 3'd0;
    assign memory3b[336 ] = 3'd6;
    assign memory3b[337 ] = 3'd6;
    assign memory3b[338 ] = 3'd0;
    assign memory3b[339 ] = 3'd6;
    assign memory3b[340 ] = 3'd6;
    assign memory3b[341 ] = 3'd6;
    assign memory3b[342 ] = 3'd0;
    assign memory3b[343 ] = 3'd1;
    assign memory3b[344 ] = 3'd1;
    assign memory3b[345 ] = 3'd2;
    assign memory3b[346 ] = 3'd0;
    assign memory3b[347 ] = 3'd0;
    assign memory3b[348 ] = 3'd0;
    assign memory3b[349 ] = 3'd0;
    assign memory3b[350 ] = 3'd2;
    assign memory3b[351 ] = 3'd0;
    assign memory3b[352 ] = 3'd0;
    assign memory3b[353 ] = 3'd0;
    assign memory3b[354 ] = 3'd0;
    assign memory3b[355 ] = 3'd3;
    assign memory3b[356 ] = 3'd2;
    assign memory3b[357 ] = 3'd0;
    assign memory3b[358 ] = 3'd0;
    assign memory3b[359 ] = 3'd0;
    assign memory3b[360 ] = 3'd3;
    assign memory3b[361 ] = 3'd3;
    assign memory3b[362 ] = 3'd0;
    assign memory3b[363 ] = 3'd0;
    assign memory3b[364 ] = 3'd0;
    assign memory3b[365 ] = 3'd0;
    assign memory3b[366 ] = 3'd0;
    assign memory3b[367 ] = 3'd3;
    assign memory3b[368 ] = 3'd6;
    assign memory3b[369 ] = 3'd6;
    assign memory3b[370 ] = 3'd6;
    assign memory3b[371 ] = 3'd6;
    assign memory3b[372 ] = 3'd6;
    assign memory3b[373 ] = 3'd6;
    assign memory3b[374 ] = 3'd2;
    assign memory3b[375 ] = 3'd0;
    assign memory3b[376 ] = 3'd2;
    assign memory3b[377 ] = 3'd3;
    assign memory3b[378 ] = 3'd3;
    assign memory3b[379 ] = 3'd0;
    assign memory3b[380 ] = 3'd1;
    assign memory3b[381 ] = 3'd0;
    assign memory3b[382 ] = 3'd3;
    assign memory3b[383 ] = 3'd0;
    assign memory3b[384 ] = 3'd3;
    assign memory3b[385 ] = 3'd3;
    assign memory3b[386 ] = 3'd0;
    assign memory3b[387 ] = 3'd0;
    assign memory3b[388 ] = 3'd2;
    assign memory3b[389 ] = 3'd2;
    assign memory3b[390 ] = 3'd2;
    assign memory3b[391 ] = 3'd0;
    assign memory3b[392 ] = 3'd0;
    assign memory3b[393 ] = 3'd0;
    assign memory3b[394 ] = 3'd1;
    assign memory3b[395 ] = 3'd0;
    assign memory3b[396 ] = 3'd0;
    assign memory3b[397 ] = 3'd0;
    assign memory3b[398 ] = 3'd0;
    assign memory3b[399 ] = 3'd0;
    assign memory3b[400 ] = 3'd3;
    assign memory3b[401 ] = 3'd3;
    assign memory3b[402 ] = 3'd0;
    assign memory3b[403 ] = 3'd3;
    assign memory3b[404 ] = 3'd0;
    assign memory3b[405 ] = 3'd3;
    assign memory3b[406 ] = 3'd3;
    assign memory3b[407 ] = 3'd0;
    assign memory3b[408 ] = 3'd0;
    assign memory3b[409 ] = 3'd0;
    assign memory3b[410 ] = 3'd0;
    assign memory3b[411 ] = 3'd1;
    assign memory3b[412 ] = 3'd1;
    assign memory3b[413 ] = 3'd0;
    assign memory3b[414 ] = 3'd0;
    assign memory3b[415 ] = 3'd0;
    assign memory3b[416 ] = 3'd0;
    assign memory3b[417 ] = 3'd0;
    assign memory3b[418 ] = 3'd0;
    assign memory3b[419 ] = 3'd0;
    assign memory3b[420 ] = 3'd0;
    assign memory3b[421 ] = 3'd0;
    assign memory3b[422 ] = 3'd3;
    assign memory3b[423 ] = 3'd3;
    assign memory3b[424 ] = 3'd0;
    assign memory3b[425 ] = 3'd0;
    assign memory3b[426 ] = 3'd0;
    assign memory3b[427 ] = 3'd0;
    assign memory3b[428 ] = 3'd0;
    assign memory3b[429 ] = 3'd0;
    assign memory3b[430 ] = 3'd2;
    assign memory3b[431 ] = 3'd0;
    assign memory3b[432 ] = 3'd3;
    assign memory3b[433 ] = 3'd3;
    assign memory3b[434 ] = 3'd0;
    assign memory3b[435 ] = 3'd3;
    assign memory3b[436 ] = 3'd0;
    assign memory3b[437 ] = 3'd3;
    assign memory3b[438 ] = 3'd3;
    assign memory3b[439 ] = 3'd0;
    assign memory3b[440 ] = 3'd0;
    assign memory3b[441 ] = 3'd0;
    assign memory3b[442 ] = 3'd0;
    assign memory3b[443 ] = 3'd0;
    assign memory3b[444 ] = 3'd0;
    assign memory3b[445 ] = 3'd0;
    assign memory3b[446 ] = 3'd0;
    assign memory3b[447 ] = 3'd1;
    assign memory3b[448 ] = 3'd0;
    assign memory3b[449 ] = 3'd0;
    assign memory3b[450 ] = 3'd0;
    assign memory3b[451 ] = 3'd0;
    assign memory3b[452 ] = 3'd0;
    assign memory3b[453 ] = 3'd0;
    assign memory3b[454 ] = 3'd0;
    assign memory3b[455 ] = 3'd0;
    assign memory3b[456 ] = 3'd0;
    assign memory3b[457 ] = 3'd0;
    assign memory3b[458 ] = 3'd0;
    assign memory3b[459 ] = 3'd0;
    assign memory3b[460 ] = 3'd0;
    assign memory3b[461 ] = 3'd0;
    assign memory3b[462 ] = 3'd0;
    assign memory3b[463 ] = 3'd1;
    assign memory3b[464 ] = 3'd3;
    assign memory3b[465 ] = 3'd0;
    assign memory3b[466 ] = 3'd0;
    assign memory3b[467 ] = 3'd3;
    assign memory3b[468 ] = 3'd0;
    assign memory3b[469 ] = 3'd0;
    assign memory3b[470 ] = 3'd0;
    assign memory3b[471 ] = 3'd1;
    assign memory3b[472 ] = 3'd0;
    assign memory3b[473 ] = 3'd0;
    assign memory3b[474 ] = 3'd1;
    assign memory3b[475 ] = 3'd0;
    assign memory3b[476 ] = 3'd0;
    assign memory3b[477 ] = 3'd0;
    assign memory3b[478 ] = 3'd0;
    assign memory3b[479 ] = 3'd0;
    assign memory3b[480 ] = 3'd0;
    assign memory3b[481 ] = 3'd0;
    assign memory3b[482 ] = 3'd0;
    assign memory3b[483 ] = 3'd0;
    assign memory3b[484 ] = 3'd0;
    assign memory3b[485 ] = 3'd0;
    assign memory3b[486 ] = 3'd3;
    assign memory3b[487 ] = 3'd0;
    assign memory3b[488 ] = 3'd0;
    assign memory3b[489 ] = 3'd0;
    assign memory3b[490 ] = 3'd0;
    assign memory3b[491 ] = 3'd0;
    assign memory3b[492 ] = 3'd0;
    assign memory3b[493 ] = 3'd2;
    assign memory3b[494 ] = 3'd0;
    assign memory3b[495 ] = 3'd0;
    assign memory3b[496 ] = 3'd0;
    assign memory3b[497 ] = 3'd0;
    assign memory3b[498 ] = 3'd2;
    assign memory3b[499 ] = 3'd0;
    assign memory3b[500 ] = 3'd0;
    assign memory3b[501 ] = 3'd0;
    assign memory3b[502 ] = 3'd0;
    assign memory3b[503 ] = 3'd3;
    assign memory3b[504 ] = 3'd1;
    assign memory3b[505 ] = 3'd0;
    assign memory3b[506 ] = 3'd3;
    assign memory3b[507 ] = 3'd0;
    assign memory3b[508 ] = 3'd0;
    assign memory3b[509 ] = 3'd0;
    assign memory3b[510 ] = 3'd1;
    assign memory3b[511 ] = 3'd0;
    assign memory3b[512 ] = 3'd0;
    assign memory3b[513 ] = 3'd0;
    assign memory3b[514 ] = 3'd0;
    assign memory3b[515 ] = 3'd0;
    assign memory3b[516 ] = 3'd0;
    assign memory3b[517 ] = 3'd3;
    assign memory3b[518 ] = 3'd0;
    assign memory3b[519 ] = 3'd0;
    assign memory3b[520 ] = 3'd1;
    assign memory3b[521 ] = 3'd0;
    assign memory3b[522 ] = 3'd1;
    assign memory3b[523 ] = 3'd0;
    assign memory3b[524 ] = 3'd0;
    assign memory3b[525 ] = 3'd1;
    assign memory3b[526 ] = 3'd0;
    assign memory3b[527 ] = 3'd0;
    assign memory3b[528 ] = 3'd0;
    assign memory3b[529 ] = 3'd0;
    assign memory3b[530 ] = 3'd0;
    assign memory3b[531 ] = 3'd0;
    assign memory3b[532 ] = 3'd0;
    assign memory3b[533 ] = 3'd0;
    assign memory3b[534 ] = 3'd0;
    assign memory3b[535 ] = 3'd1;
    assign memory3b[536 ] = 3'd3;
    assign memory3b[537 ] = 3'd0;
    assign memory3b[538 ] = 3'd0;
    assign memory3b[539 ] = 3'd2;
    assign memory3b[540 ] = 3'd0;
    assign memory3b[541 ] = 3'd0;
    assign memory3b[542 ] = 3'd0;
    assign memory3b[543 ] = 3'd3;
    assign memory3b[544 ] = 3'd1;
    assign memory3b[545 ] = 3'd0;
    assign memory3b[546 ] = 3'd0;
    assign memory3b[547 ] = 3'd0;
    assign memory3b[548 ] = 3'd0;
    assign memory3b[549 ] = 3'd0;
    assign memory3b[550 ] = 3'd0;
    assign memory3b[551 ] = 3'd0;
    assign memory3b[552 ] = 3'd0;
    assign memory3b[553 ] = 3'd0;
    assign memory3b[554 ] = 3'd0;
    assign memory3b[555 ] = 3'd1;
    assign memory3b[556 ] = 3'd0;
    assign memory3b[557 ] = 3'd0;
    assign memory3b[558 ] = 3'd1;
    assign memory3b[559 ] = 3'd0;
    assign memory3b[560 ] = 3'd0;
    assign memory3b[561 ] = 3'd1;
    assign memory3b[562 ] = 3'd1;
    assign memory3b[563 ] = 3'd1;
    assign memory3b[564 ] = 3'd0;
    assign memory3b[565 ] = 3'd0;
    assign memory3b[566 ] = 3'd0;
    assign memory3b[567 ] = 3'd0;
    assign memory3b[568 ] = 3'd1;
    assign memory3b[569 ] = 3'd0;
    assign memory3b[570 ] = 3'd0;
    assign memory3b[571 ] = 3'd0;
    assign memory3b[572 ] = 3'd0;
    assign memory3b[573 ] = 3'd0;
    assign memory3b[574 ] = 3'd0;
    assign memory3b[575 ] = 3'd0;
    assign memory3b[576 ] = 3'd0;
    assign memory3b[577 ] = 3'd0;
    assign memory3b[578 ] = 3'd0;
    assign memory3b[579 ] = 3'd0;
    assign memory3b[580 ] = 3'd0;
    assign memory3b[581 ] = 3'd0;
    assign memory3b[582 ] = 3'd1;
    assign memory3b[583 ] = 3'd0;
    assign memory3b[584 ] = 3'd0;
    assign memory3b[585 ] = 3'd0;
    assign memory3b[586 ] = 3'd0;
    assign memory3b[587 ] = 3'd0;
    assign memory3b[588 ] = 3'd0;
    assign memory3b[589 ] = 3'd0;
    assign memory3b[590 ] = 3'd0;
    assign memory3b[591 ] = 3'd0;
    assign memory3b[592 ] = 3'd0;
    assign memory3b[593 ] = 3'd0;
    assign memory3b[594 ] = 3'd0;
    assign memory3b[595 ] = 3'd3;
    assign memory3b[596 ] = 3'd0;
    assign memory3b[597 ] = 3'd0;
    assign memory3b[598 ] = 3'd0;
    assign memory3b[599 ] = 3'd1;
    assign memory3b[600 ] = 3'd3;
    assign memory3b[601 ] = 3'd0;
    assign memory3b[602 ] = 3'd0;
    assign memory3b[603 ] = 3'd0;
    assign memory3b[604 ] = 3'd0;
    assign memory3b[605 ] = 3'd0;
    assign memory3b[606 ] = 3'd3;
    assign memory3b[607 ] = 3'd0;
    assign memory3b[608 ] = 3'd3;
    assign memory3b[609 ] = 3'd3;
    assign memory3b[610 ] = 3'd0;
    assign memory3b[611 ] = 3'd0;
    assign memory3b[612 ] = 3'd0;
    assign memory3b[613 ] = 3'd0;
    assign memory3b[614 ] = 3'd0;
    assign memory3b[615 ] = 3'd0;
    assign memory3b[616 ] = 3'd0;
    assign memory3b[617 ] = 3'd0;
    assign memory3b[618 ] = 3'd0;
    assign memory3b[619 ] = 3'd0;
    assign memory3b[620 ] = 3'd1;
    assign memory3b[621 ] = 3'd3;
    assign memory3b[622 ] = 3'd0;
    assign memory3b[623 ] = 3'd0;
    assign memory3b[624 ] = 3'd1;
    assign memory3b[625 ] = 3'd0;
    assign memory3b[626 ] = 3'd1;
    assign memory3b[627 ] = 3'd0;
    assign memory3b[628 ] = 3'd0;
    assign memory3b[629 ] = 3'd3;
    assign memory3b[630 ] = 3'd0;
    assign memory3b[631 ] = 3'd3;
    assign memory3b[632 ] = 3'd0;
    assign memory3b[633 ] = 3'd0;
    assign memory3b[634 ] = 3'd0;
    assign memory3b[635 ] = 3'd3;
    assign memory3b[636 ] = 3'd0;
    assign memory3b[637 ] = 3'd0;
    assign memory3b[638 ] = 3'd0;
    assign memory3b[639 ] = 3'd0;
    assign memory3b[640 ] = 3'd0;
    assign memory3b[641 ] = 3'd0;
    assign memory3b[642 ] = 3'd0;
    assign memory3b[643 ] = 3'd0;
    assign memory3b[644 ] = 3'd0;
    assign memory3b[645 ] = 3'd0;
    assign memory3b[646 ] = 3'd0;
    assign memory3b[647 ] = 3'd0;
    assign memory3b[648 ] = 3'd0;
    assign memory3b[649 ] = 3'd0;
    assign memory3b[650 ] = 3'd0;
    assign memory3b[651 ] = 3'd0;
    assign memory3b[652 ] = 3'd0;
    assign memory3b[653 ] = 3'd0;
    assign memory3b[654 ] = 3'd0;
    assign memory3b[655 ] = 3'd0;
    assign memory3b[656 ] = 3'd3;
    assign memory3b[657 ] = 3'd0;
    assign memory3b[658 ] = 3'd0;
    assign memory3b[659 ] = 3'd0;
    assign memory3b[660 ] = 3'd0;
    assign memory3b[661 ] = 3'd0;
    assign memory3b[662 ] = 3'd0;
    assign memory3b[663 ] = 3'd0;
    assign memory3b[664 ] = 3'd0;
    assign memory3b[665 ] = 3'd0;
    assign memory3b[666 ] = 3'd0;
    assign memory3b[667 ] = 3'd0;
    assign memory3b[668 ] = 3'd0;
    assign memory3b[669 ] = 3'd0;
    assign memory3b[670 ] = 3'd0;
    assign memory3b[671 ] = 3'd0;
    assign memory3b[672 ] = 3'd3;
    assign memory3b[673 ] = 3'd0;
    assign memory3b[674 ] = 3'd0;
    assign memory3b[675 ] = 3'd0;
    assign memory3b[676 ] = 3'd0;
    assign memory3b[677 ] = 3'd0;
    assign memory3b[678 ] = 3'd0;
    assign memory3b[679 ] = 3'd4;
    assign memory3b[680 ] = 3'd5;
    assign memory3b[681 ] = 3'd0;
    assign memory3b[682 ] = 3'd0;
    assign memory3b[683 ] = 3'd0;
    assign memory3b[684 ] = 3'd0;
    assign memory3b[685 ] = 3'd0;
    assign memory3b[686 ] = 3'd0;
    assign memory3b[687 ] = 3'd0;
    assign memory3b[688 ] = 3'd0;
    assign memory3b[689 ] = 3'd0;
    assign memory3b[690 ] = 3'd0;
    assign memory3b[691 ] = 3'd0;
    assign memory3b[692 ] = 3'd0;
    assign memory3b[693 ] = 3'd0;
    assign memory3b[694 ] = 3'd0;
    assign memory3b[695 ] = 3'd0;
    assign memory3b[696 ] = 3'd0;
    assign memory3b[697 ] = 3'd0;
    assign memory3b[698 ] = 3'd0;
    assign memory3b[699 ] = 3'd0;
    assign memory3b[700 ] = 3'd0;
    assign memory3b[701 ] = 3'd0;
    assign memory3b[702 ] = 3'd0;
    assign memory3b[703 ] = 3'd0;
    assign memory3b[704 ] = 3'd0;
    assign memory3b[705 ] = 3'd0;
    assign memory3b[706 ] = 3'd0;
    assign memory3b[707 ] = 3'd0;
    assign memory3b[708 ] = 3'd0;
    assign memory3b[709 ] = 3'd0;
    assign memory3b[710 ] = 3'd4;
    assign memory3b[711 ] = 3'd4;
    assign memory3b[712 ] = 3'd5;
    assign memory3b[713 ] = 3'd5;
    assign memory3b[714 ] = 3'd1;
    assign memory3b[715 ] = 3'd0;
    assign memory3b[716 ] = 3'd0;
    assign memory3b[717 ] = 3'd0;
    assign memory3b[718 ] = 3'd0;
    assign memory3b[719 ] = 3'd0;
    assign memory3b[720 ] = 3'd3;
    assign memory3b[721 ] = 3'd0;
    assign memory3b[722 ] = 3'd0;
    assign memory3b[723 ] = 3'd1;
    assign memory3b[724 ] = 3'd0;
    assign memory3b[725 ] = 3'd0;
    assign memory3b[726 ] = 3'd0;
    assign memory3b[727 ] = 3'd0;
    assign memory3b[728 ] = 3'd0;
    assign memory3b[729 ] = 3'd0;
    assign memory3b[730 ] = 3'd0;
    assign memory3b[731 ] = 3'd0;
    assign memory3b[732 ] = 3'd0;
    assign memory3b[733 ] = 3'd0;
    assign memory3b[734 ] = 3'd0;
    assign memory3b[735 ] = 3'd0;
    assign memory3b[736 ] = 3'd0;
    assign memory3b[737 ] = 3'd0;
    assign memory3b[738 ] = 3'd0;
    assign memory3b[739 ] = 3'd0;
    assign memory3b[740 ] = 3'd0;
    assign memory3b[741 ] = 3'd4;
    assign memory3b[742 ] = 3'd4;
    assign memory3b[743 ] = 3'd4;
    assign memory3b[744 ] = 3'd4;
    assign memory3b[745 ] = 3'd5;
    assign memory3b[746 ] = 3'd5;
    assign memory3b[747 ] = 3'd3;
    assign memory3b[748 ] = 3'd0;
    assign memory3b[749 ] = 3'd0;
    assign memory3b[750 ] = 3'd0;
    assign memory3b[751 ] = 3'd6;
    assign memory3b[752 ] = 3'd0;
    assign memory3b[753 ] = 3'd6;
    assign memory3b[754 ] = 3'd0;
    assign memory3b[755 ] = 3'd0;
    assign memory3b[756 ] = 3'd0;
    assign memory3b[757 ] = 3'd0;
    assign memory3b[758 ] = 3'd0;
    assign memory3b[759 ] = 3'd0;
    assign memory3b[760 ] = 3'd0;
    assign memory3b[761 ] = 3'd0;
    assign memory3b[762 ] = 3'd0;
    assign memory3b[763 ] = 3'd0;
    assign memory3b[764 ] = 3'd0;
    assign memory3b[765 ] = 3'd0;
    assign memory3b[766 ] = 3'd0;
    assign memory3b[767 ] = 3'd0;
    assign memory3b[768 ] = 3'd0;
    assign memory3b[769 ] = 3'd0;
    assign memory3b[770 ] = 3'd0;
    assign memory3b[771 ] = 3'd0;
    assign memory3b[772 ] = 3'd1;
    assign memory3b[773 ] = 3'd4;
    assign memory3b[774 ] = 3'd4;
    assign memory3b[775 ] = 3'd4;
    assign memory3b[776 ] = 3'd4;
    assign memory3b[777 ] = 3'd5;
    assign memory3b[778 ] = 3'd1;
    assign memory3b[779 ] = 3'd0;
    assign memory3b[780 ] = 3'd0;
    assign memory3b[781 ] = 3'd6;
    assign memory3b[782 ] = 3'd6;
    assign memory3b[783 ] = 3'd6;
    assign memory3b[784 ] = 3'd6;
    assign memory3b[785 ] = 3'd6;
    assign memory3b[786 ] = 3'd6;
    assign memory3b[787 ] = 3'd0;
    assign memory3b[788 ] = 3'd0;
    assign memory3b[789 ] = 3'd0;
    assign memory3b[790 ] = 3'd1;
    assign memory3b[791 ] = 3'd0;
    assign memory3b[792 ] = 3'd0;
    assign memory3b[793 ] = 3'd0;
    assign memory3b[794 ] = 3'd0;
    assign memory3b[795 ] = 3'd3;
    assign memory3b[796 ] = 3'd0;
    assign memory3b[797 ] = 3'd0;
    assign memory3b[798 ] = 3'd0;
    assign memory3b[799 ] = 3'd0;
    assign memory3b[800 ] = 3'd0;
    assign memory3b[801 ] = 3'd0;
    assign memory3b[802 ] = 3'd0;
    assign memory3b[803 ] = 3'd0;
    assign memory3b[804 ] = 3'd0;
    assign memory3b[805 ] = 3'd0;
    assign memory3b[806 ] = 3'd2;
    assign memory3b[807 ] = 3'd3;
    assign memory3b[808 ] = 3'd0;
    assign memory3b[809 ] = 3'd0;
    assign memory3b[810 ] = 3'd1;
    assign memory3b[811 ] = 3'd1;
    assign memory3b[812 ] = 3'd2;
    assign memory3b[813 ] = 3'd0;
    assign memory3b[814 ] = 3'd3;
    assign memory3b[815 ] = 3'd3;
    assign memory3b[816 ] = 3'd0;
    assign memory3b[817 ] = 3'd0;
    assign memory3b[818 ] = 3'd0;
    assign memory3b[819 ] = 3'd0;
    assign memory3b[820 ] = 3'd1;
    assign memory3b[821 ] = 3'd2;
    assign memory3b[822 ] = 3'd0;
    assign memory3b[823 ] = 3'd0;
    assign memory3b[824 ] = 3'd0;
    assign memory3b[825 ] = 3'd0;
    assign memory3b[826 ] = 3'd0;
    assign memory3b[827 ] = 3'd0;
    assign memory3b[828 ] = 3'd0;
    assign memory3b[829 ] = 3'd0;
    assign memory3b[830 ] = 3'd0;
    assign memory3b[831 ] = 3'd0;
    assign memory3b[832 ] = 3'd0;
    assign memory3b[833 ] = 3'd0;
    assign memory3b[834 ] = 3'd0;
    assign memory3b[835 ] = 3'd3;
    assign memory3b[836 ] = 3'd1;
    assign memory3b[837 ] = 3'd0;
    assign memory3b[838 ] = 3'd0;
    assign memory3b[839 ] = 3'd3;
    assign memory3b[840 ] = 3'd0;
    assign memory3b[841 ] = 3'd0;
    assign memory3b[842 ] = 3'd0;
    assign memory3b[843 ] = 3'd0;
    assign memory3b[844 ] = 3'd0;
    assign memory3b[845 ] = 3'd0;
    assign memory3b[846 ] = 3'd0;
    assign memory3b[847 ] = 3'd0;
    assign memory3b[848 ] = 3'd0;
    assign memory3b[849 ] = 3'd0;
    assign memory3b[850 ] = 3'd3;
    assign memory3b[851 ] = 3'd0;
    assign memory3b[852 ] = 3'd3;
    assign memory3b[853 ] = 3'd0;
    assign memory3b[854 ] = 3'd0;
    assign memory3b[855 ] = 3'd0;
    assign memory3b[856 ] = 3'd0;
    assign memory3b[857 ] = 3'd0;
    assign memory3b[858 ] = 3'd0;
    assign memory3b[859 ] = 3'd1;
    assign memory3b[860 ] = 3'd0;
    assign memory3b[861 ] = 3'd0;
    assign memory3b[862 ] = 3'd0;
    assign memory3b[863 ] = 3'd0;
    assign memory3b[864 ] = 3'd0;
    assign memory3b[865 ] = 3'd0;
    assign memory3b[866 ] = 3'd0;
    assign memory3b[867 ] = 3'd0;
    assign memory3b[868 ] = 3'd0;
    assign memory3b[869 ] = 3'd2;
    assign memory3b[870 ] = 3'd0;
    assign memory3b[871 ] = 3'd0;
    assign memory3b[872 ] = 3'd0;
    assign memory3b[873 ] = 3'd2;
    assign memory3b[874 ] = 3'd0;
    assign memory3b[875 ] = 3'd0;
    assign memory3b[876 ] = 3'd3;
    assign memory3b[877 ] = 3'd3;
    assign memory3b[878 ] = 3'd0;
    assign memory3b[879 ] = 3'd0;
    assign memory3b[880 ] = 3'd0;
    assign memory3b[881 ] = 3'd0;
    assign memory3b[882 ] = 3'd0;
    assign memory3b[883 ] = 3'd0;
    assign memory3b[884 ] = 3'd0;
    assign memory3b[885 ] = 3'd1;
    assign memory3b[886 ] = 3'd0;
    assign memory3b[887 ] = 3'd0;
    assign memory3b[888 ] = 3'd0;
    assign memory3b[889 ] = 3'd0;
    assign memory3b[890 ] = 3'd0;
    assign memory3b[891 ] = 3'd0;
    assign memory3b[892 ] = 3'd3;
    assign memory3b[893 ] = 3'd0;
    assign memory3b[894 ] = 3'd2;
    assign memory3b[895 ] = 3'd0;
    assign memory3b[896 ] = 3'd0;
    assign memory3b[897 ] = 3'd3;
    assign memory3b[898 ] = 3'd0;
    assign memory3b[899 ] = 3'd3;
    assign memory3b[900 ] = 3'd0;
    assign memory3b[901 ] = 3'd0;
    assign memory3b[902 ] = 3'd0;
    assign memory3b[903 ] = 3'd0;
    assign memory3b[904 ] = 3'd0;
    assign memory3b[905 ] = 3'd0;
    assign memory3b[906 ] = 3'd0;
    assign memory3b[907 ] = 3'd2;
    assign memory3b[908 ] = 3'd2;
    assign memory3b[909 ] = 3'd0;
    assign memory3b[910 ] = 3'd0;
    assign memory3b[911 ] = 3'd0;
    assign memory3b[912 ] = 3'd0;
    assign memory3b[913 ] = 3'd3;
    assign memory3b[914 ] = 3'd0;
    assign memory3b[915 ] = 3'd0;
    assign memory3b[916 ] = 3'd0;
    assign memory3b[917 ] = 3'd0;
    assign memory3b[918 ] = 3'd0;
    assign memory3b[919 ] = 3'd0;
    assign memory3b[920 ] = 3'd0;
    assign memory3b[921 ] = 3'd0;
    assign memory3b[922 ] = 3'd0;
    assign memory3b[923 ] = 3'd0;
    assign memory3b[924 ] = 3'd0;
    assign memory3b[925 ] = 3'd0;
    assign memory3b[926 ] = 3'd0;
    assign memory3b[927 ] = 3'd1;
    assign memory3b[928 ] = 3'd0;
    assign memory3b[929 ] = 3'd0;
    assign memory3b[930 ] = 3'd0;
    assign memory3b[931 ] = 3'd0;
    assign memory3b[932 ] = 3'd0;
    assign memory3b[933 ] = 3'd0;
    assign memory3b[934 ] = 3'd1;
    assign memory3b[935 ] = 3'd0;
    assign memory3b[936 ] = 3'd3;
    assign memory3b[937 ] = 3'd0;
    assign memory3b[938 ] = 3'd0;
    assign memory3b[939 ] = 3'd0;
    assign memory3b[940 ] = 3'd0;
    assign memory3b[941 ] = 3'd0;
    assign memory3b[942 ] = 3'd0;
    assign memory3b[943 ] = 3'd0;
    assign memory3b[944 ] = 3'd0;
    assign memory3b[945 ] = 3'd0;
    assign memory3b[946 ] = 3'd0;
    assign memory3b[947 ] = 3'd0;
    assign memory3b[948 ] = 3'd0;
    assign memory3b[949 ] = 3'd0;
    assign memory3b[950 ] = 3'd0;
    assign memory3b[951 ] = 3'd0;
    assign memory3b[952 ] = 3'd0;
    assign memory3b[953 ] = 3'd0;
    assign memory3b[954 ] = 3'd0;
    assign memory3b[955 ] = 3'd0;
    assign memory3b[956 ] = 3'd0;
    assign memory3b[957 ] = 3'd0;
    assign memory3b[958 ] = 3'd0;
    assign memory3b[959 ] = 3'd3;
    assign memory3b[960 ] = 3'd0;
    assign memory3b[961 ] = 3'd0;
    assign memory3b[962 ] = 3'd0;
    assign memory3b[963 ] = 3'd0;
    assign memory3b[964 ] = 3'd0;
    assign memory3b[965 ] = 3'd0;
    assign memory3b[966 ] = 3'd0;
    assign memory3b[967 ] = 3'd0;
    assign memory3b[968 ] = 3'd0;
    assign memory3b[969 ] = 3'd3;
    assign memory3b[970 ] = 3'd0;
    assign memory3b[971 ] = 3'd0;
    assign memory3b[972 ] = 3'd0;
    assign memory3b[973 ] = 3'd3;
    assign memory3b[974 ] = 3'd1;
    assign memory3b[975 ] = 3'd3;
    assign memory3b[976 ] = 3'd0;
    assign memory3b[977 ] = 3'd0;
    assign memory3b[978 ] = 3'd0;
    assign memory3b[979 ] = 3'd1;
    assign memory3b[980 ] = 3'd0;
    assign memory3b[981 ] = 3'd0;
    assign memory3b[982 ] = 3'd0;
    assign memory3b[983 ] = 3'd0;
    assign memory3b[984 ] = 3'd3;
    assign memory3b[985 ] = 3'd2;
    assign memory3b[986 ] = 3'd0;
    assign memory3b[987 ] = 3'd1;
    assign memory3b[988 ] = 3'd0;
    assign memory3b[989 ] = 3'd0;
    assign memory3b[990 ] = 3'd0;
    assign memory3b[991 ] = 3'd0;
    assign memory3b[992 ] = 3'd0;
    assign memory3b[993 ] = 3'd0;
    assign memory3b[994 ] = 3'd0;
    assign memory3b[995 ] = 3'd0;
    assign memory3b[996 ] = 3'd0;
    assign memory3b[997 ] = 3'd0;
    assign memory3b[998 ] = 3'd0;
    assign memory3b[999 ] = 3'd0;
    assign memory3b[1000] = 3'd0;
    assign memory3b[1001] = 3'd0;
    assign memory3b[1002] = 3'd0;
    assign memory3b[1003] = 3'd0;
    assign memory3b[1004] = 3'd1;
    assign memory3b[1005] = 3'd0;
    assign memory3b[1006] = 3'd3;
    assign memory3b[1007] = 3'd0;
    assign memory3b[1008] = 3'd0;
    assign memory3b[1009] = 3'd0;
    assign memory3b[1010] = 3'd0;
    assign memory3b[1011] = 3'd0;
    assign memory3b[1012] = 3'd0;
    assign memory3b[1013] = 3'd0;
    assign memory3b[1014] = 3'd0;
    assign memory3b[1015] = 3'd0;
    assign memory3b[1016] = 3'd0;
    assign memory3b[1017] = 3'd0;
    assign memory3b[1018] = 3'd2;
    assign memory3b[1019] = 3'd0;
    assign memory3b[1020] = 3'd0;
    assign memory3b[1021] = 3'd0;
    assign memory3b[1022] = 3'd0;
    assign memory3b[1023] = 3'd0;

    assign memory4a[0   ] = 3'd0;
    assign memory4a[1   ] = 3'd1;
    assign memory4a[2   ] = 3'd2;
    assign memory4a[3   ] = 3'd2;
    assign memory4a[4   ] = 3'd2;
    assign memory4a[5   ] = 3'd2;
    assign memory4a[6   ] = 3'd2;
    assign memory4a[7   ] = 3'd2;
    assign memory4a[8   ] = 3'd2;
    assign memory4a[9   ] = 3'd2;
    assign memory4a[10  ] = 3'd2;
    assign memory4a[11  ] = 3'd2;
    assign memory4a[12  ] = 3'd2;
    assign memory4a[13  ] = 3'd2;
    assign memory4a[14  ] = 3'd2;
    assign memory4a[15  ] = 3'd2;
    assign memory4a[16  ] = 3'd2;
    assign memory4a[17  ] = 3'd2;
    assign memory4a[18  ] = 3'd2;
    assign memory4a[19  ] = 3'd2;
    assign memory4a[20  ] = 3'd2;
    assign memory4a[21  ] = 3'd2;
    assign memory4a[22  ] = 3'd2;
    assign memory4a[23  ] = 3'd2;
    assign memory4a[24  ] = 3'd2;
    assign memory4a[25  ] = 3'd2;
    assign memory4a[26  ] = 3'd2;
    assign memory4a[27  ] = 3'd2;
    assign memory4a[28  ] = 3'd2;
    assign memory4a[29  ] = 3'd2;
    assign memory4a[30  ] = 3'd1;
    assign memory4a[31  ] = 3'd0;
    assign memory4a[32  ] = 3'd1;
    assign memory4a[33  ] = 3'd0;
    assign memory4a[34  ] = 3'd1;
    assign memory4a[35  ] = 3'd2;
    assign memory4a[36  ] = 3'd2;
    assign memory4a[37  ] = 3'd2;
    assign memory4a[38  ] = 3'd2;
    assign memory4a[39  ] = 3'd2;
    assign memory4a[40  ] = 3'd2;
    assign memory4a[41  ] = 3'd2;
    assign memory4a[42  ] = 3'd2;
    assign memory4a[43  ] = 3'd2;
    assign memory4a[44  ] = 3'd2;
    assign memory4a[45  ] = 3'd2;
    assign memory4a[46  ] = 3'd2;
    assign memory4a[47  ] = 3'd2;
    assign memory4a[48  ] = 3'd2;
    assign memory4a[49  ] = 3'd2;
    assign memory4a[50  ] = 3'd2;
    assign memory4a[51  ] = 3'd2;
    assign memory4a[52  ] = 3'd2;
    assign memory4a[53  ] = 3'd2;
    assign memory4a[54  ] = 3'd2;
    assign memory4a[55  ] = 3'd2;
    assign memory4a[56  ] = 3'd2;
    assign memory4a[57  ] = 3'd2;
    assign memory4a[58  ] = 3'd2;
    assign memory4a[59  ] = 3'd2;
    assign memory4a[60  ] = 3'd2;
    assign memory4a[61  ] = 3'd1;
    assign memory4a[62  ] = 3'd0;
    assign memory4a[63  ] = 3'd1;
    assign memory4a[64  ] = 3'd2;
    assign memory4a[65  ] = 3'd1;
    assign memory4a[66  ] = 3'd0;
    assign memory4a[67  ] = 3'd1;
    assign memory4a[68  ] = 3'd2;
    assign memory4a[69  ] = 3'd2;
    assign memory4a[70  ] = 3'd2;
    assign memory4a[71  ] = 3'd2;
    assign memory4a[72  ] = 3'd2;
    assign memory4a[73  ] = 3'd2;
    assign memory4a[74  ] = 3'd2;
    assign memory4a[75  ] = 3'd2;
    assign memory4a[76  ] = 3'd2;
    assign memory4a[77  ] = 3'd2;
    assign memory4a[78  ] = 3'd2;
    assign memory4a[79  ] = 3'd2;
    assign memory4a[80  ] = 3'd2;
    assign memory4a[81  ] = 3'd2;
    assign memory4a[82  ] = 3'd2;
    assign memory4a[83  ] = 3'd2;
    assign memory4a[84  ] = 3'd2;
    assign memory4a[85  ] = 3'd2;
    assign memory4a[86  ] = 3'd2;
    assign memory4a[87  ] = 3'd2;
    assign memory4a[88  ] = 3'd2;
    assign memory4a[89  ] = 3'd2;
    assign memory4a[90  ] = 3'd2;
    assign memory4a[91  ] = 3'd2;
    assign memory4a[92  ] = 3'd1;
    assign memory4a[93  ] = 3'd0;
    assign memory4a[94  ] = 3'd1;
    assign memory4a[95  ] = 3'd2;
    assign memory4a[96  ] = 3'd2;
    assign memory4a[97  ] = 3'd2;
    assign memory4a[98  ] = 3'd1;
    assign memory4a[99  ] = 3'd0;
    assign memory4a[100 ] = 3'd1;
    assign memory4a[101 ] = 3'd2;
    assign memory4a[102 ] = 3'd2;
    assign memory4a[103 ] = 3'd2;
    assign memory4a[104 ] = 3'd2;
    assign memory4a[105 ] = 3'd2;
    assign memory4a[106 ] = 3'd2;
    assign memory4a[107 ] = 3'd2;
    assign memory4a[108 ] = 3'd2;
    assign memory4a[109 ] = 3'd2;
    assign memory4a[110 ] = 3'd2;
    assign memory4a[111 ] = 3'd2;
    assign memory4a[112 ] = 3'd2;
    assign memory4a[113 ] = 3'd2;
    assign memory4a[114 ] = 3'd2;
    assign memory4a[115 ] = 3'd2;
    assign memory4a[116 ] = 3'd2;
    assign memory4a[117 ] = 3'd2;
    assign memory4a[118 ] = 3'd2;
    assign memory4a[119 ] = 3'd2;
    assign memory4a[120 ] = 3'd2;
    assign memory4a[121 ] = 3'd2;
    assign memory4a[122 ] = 3'd2;
    assign memory4a[123 ] = 3'd1;
    assign memory4a[124 ] = 3'd0;
    assign memory4a[125 ] = 3'd1;
    assign memory4a[126 ] = 3'd2;
    assign memory4a[127 ] = 3'd2;
    assign memory4a[128 ] = 3'd2;
    assign memory4a[129 ] = 3'd2;
    assign memory4a[130 ] = 3'd2;
    assign memory4a[131 ] = 3'd1;
    assign memory4a[132 ] = 3'd0;
    assign memory4a[133 ] = 3'd1;
    assign memory4a[134 ] = 3'd2;
    assign memory4a[135 ] = 3'd2;
    assign memory4a[136 ] = 3'd2;
    assign memory4a[137 ] = 3'd2;
    assign memory4a[138 ] = 3'd2;
    assign memory4a[139 ] = 3'd2;
    assign memory4a[140 ] = 3'd2;
    assign memory4a[141 ] = 3'd2;
    assign memory4a[142 ] = 3'd2;
    assign memory4a[143 ] = 3'd2;
    assign memory4a[144 ] = 3'd2;
    assign memory4a[145 ] = 3'd2;
    assign memory4a[146 ] = 3'd2;
    assign memory4a[147 ] = 3'd2;
    assign memory4a[148 ] = 3'd2;
    assign memory4a[149 ] = 3'd2;
    assign memory4a[150 ] = 3'd2;
    assign memory4a[151 ] = 3'd2;
    assign memory4a[152 ] = 3'd2;
    assign memory4a[153 ] = 3'd2;
    assign memory4a[154 ] = 3'd1;
    assign memory4a[155 ] = 3'd0;
    assign memory4a[156 ] = 3'd1;
    assign memory4a[157 ] = 3'd2;
    assign memory4a[158 ] = 3'd2;
    assign memory4a[159 ] = 3'd2;
    assign memory4a[160 ] = 3'd2;
    assign memory4a[161 ] = 3'd2;
    assign memory4a[162 ] = 3'd2;
    assign memory4a[163 ] = 3'd2;
    assign memory4a[164 ] = 3'd3;
    assign memory4a[165 ] = 3'd0;
    assign memory4a[166 ] = 3'd1;
    assign memory4a[167 ] = 3'd2;
    assign memory4a[168 ] = 3'd2;
    assign memory4a[169 ] = 3'd2;
    assign memory4a[170 ] = 3'd2;
    assign memory4a[171 ] = 3'd2;
    assign memory4a[172 ] = 3'd2;
    assign memory4a[173 ] = 3'd2;
    assign memory4a[174 ] = 3'd2;
    assign memory4a[175 ] = 3'd2;
    assign memory4a[176 ] = 3'd2;
    assign memory4a[177 ] = 3'd2;
    assign memory4a[178 ] = 3'd2;
    assign memory4a[179 ] = 3'd2;
    assign memory4a[180 ] = 3'd2;
    assign memory4a[181 ] = 3'd2;
    assign memory4a[182 ] = 3'd2;
    assign memory4a[183 ] = 3'd2;
    assign memory4a[184 ] = 3'd2;
    assign memory4a[185 ] = 3'd1;
    assign memory4a[186 ] = 3'd0;
    assign memory4a[187 ] = 3'd1;
    assign memory4a[188 ] = 3'd2;
    assign memory4a[189 ] = 3'd2;
    assign memory4a[190 ] = 3'd2;
    assign memory4a[191 ] = 3'd2;
    assign memory4a[192 ] = 3'd2;
    assign memory4a[193 ] = 3'd4;
    assign memory4a[194 ] = 3'd2;
    assign memory4a[195 ] = 3'd3;
    assign memory4a[196 ] = 3'd3;
    assign memory4a[197 ] = 3'd2;
    assign memory4a[198 ] = 3'd4;
    assign memory4a[199 ] = 3'd1;
    assign memory4a[200 ] = 3'd2;
    assign memory4a[201 ] = 3'd2;
    assign memory4a[202 ] = 3'd2;
    assign memory4a[203 ] = 3'd2;
    assign memory4a[204 ] = 3'd2;
    assign memory4a[205 ] = 3'd2;
    assign memory4a[206 ] = 3'd2;
    assign memory4a[207 ] = 3'd2;
    assign memory4a[208 ] = 3'd2;
    assign memory4a[209 ] = 3'd2;
    assign memory4a[210 ] = 3'd2;
    assign memory4a[211 ] = 3'd2;
    assign memory4a[212 ] = 3'd2;
    assign memory4a[213 ] = 3'd2;
    assign memory4a[214 ] = 3'd2;
    assign memory4a[215 ] = 3'd2;
    assign memory4a[216 ] = 3'd1;
    assign memory4a[217 ] = 3'd0;
    assign memory4a[218 ] = 3'd1;
    assign memory4a[219 ] = 3'd2;
    assign memory4a[220 ] = 3'd2;
    assign memory4a[221 ] = 3'd2;
    assign memory4a[222 ] = 3'd2;
    assign memory4a[223 ] = 3'd2;
    assign memory4a[224 ] = 3'd2;
    assign memory4a[225 ] = 3'd4;
    assign memory4a[226 ] = 3'd2;
    assign memory4a[227 ] = 3'd3;
    assign memory4a[228 ] = 3'd3;
    assign memory4a[229 ] = 3'd2;
    assign memory4a[230 ] = 3'd4;
    assign memory4a[231 ] = 3'd0;
    assign memory4a[232 ] = 3'd1;
    assign memory4a[233 ] = 3'd2;
    assign memory4a[234 ] = 3'd2;
    assign memory4a[235 ] = 3'd2;
    assign memory4a[236 ] = 3'd2;
    assign memory4a[237 ] = 3'd2;
    assign memory4a[238 ] = 3'd2;
    assign memory4a[239 ] = 3'd2;
    assign memory4a[240 ] = 3'd2;
    assign memory4a[241 ] = 3'd2;
    assign memory4a[242 ] = 3'd2;
    assign memory4a[243 ] = 3'd2;
    assign memory4a[244 ] = 3'd2;
    assign memory4a[245 ] = 3'd2;
    assign memory4a[246 ] = 3'd2;
    assign memory4a[247 ] = 3'd1;
    assign memory4a[248 ] = 3'd0;
    assign memory4a[249 ] = 3'd1;
    assign memory4a[250 ] = 3'd2;
    assign memory4a[251 ] = 3'd2;
    assign memory4a[252 ] = 3'd2;
    assign memory4a[253 ] = 3'd2;
    assign memory4a[254 ] = 3'd2;
    assign memory4a[255 ] = 3'd2;
    assign memory4a[256 ] = 3'd2;
    assign memory4a[257 ] = 3'd4;
    assign memory4a[258 ] = 3'd5;
    assign memory4a[259 ] = 3'd5;
    assign memory4a[260 ] = 3'd5;
    assign memory4a[261 ] = 3'd5;
    assign memory4a[262 ] = 3'd4;
    assign memory4a[263 ] = 3'd1;
    assign memory4a[264 ] = 3'd0;
    assign memory4a[265 ] = 3'd1;
    assign memory4a[266 ] = 3'd2;
    assign memory4a[267 ] = 3'd2;
    assign memory4a[268 ] = 3'd2;
    assign memory4a[269 ] = 3'd2;
    assign memory4a[270 ] = 3'd2;
    assign memory4a[271 ] = 3'd2;
    assign memory4a[272 ] = 3'd2;
    assign memory4a[273 ] = 3'd2;
    assign memory4a[274 ] = 3'd2;
    assign memory4a[275 ] = 3'd2;
    assign memory4a[276 ] = 3'd2;
    assign memory4a[277 ] = 3'd2;
    assign memory4a[278 ] = 3'd1;
    assign memory4a[279 ] = 3'd0;
    assign memory4a[280 ] = 3'd1;
    assign memory4a[281 ] = 3'd2;
    assign memory4a[282 ] = 3'd2;
    assign memory4a[283 ] = 3'd2;
    assign memory4a[284 ] = 3'd2;
    assign memory4a[285 ] = 3'd2;
    assign memory4a[286 ] = 3'd2;
    assign memory4a[287 ] = 3'd2;
    assign memory4a[288 ] = 3'd2;
    assign memory4a[289 ] = 3'd4;
    assign memory4a[290 ] = 3'd5;
    assign memory4a[291 ] = 3'd5;
    assign memory4a[292 ] = 3'd5;
    assign memory4a[293 ] = 3'd5;
    assign memory4a[294 ] = 3'd4;
    assign memory4a[295 ] = 3'd2;
    assign memory4a[296 ] = 3'd1;
    assign memory4a[297 ] = 3'd0;
    assign memory4a[298 ] = 3'd1;
    assign memory4a[299 ] = 3'd2;
    assign memory4a[300 ] = 3'd2;
    assign memory4a[301 ] = 3'd2;
    assign memory4a[302 ] = 3'd2;
    assign memory4a[303 ] = 3'd2;
    assign memory4a[304 ] = 3'd2;
    assign memory4a[305 ] = 3'd2;
    assign memory4a[306 ] = 3'd2;
    assign memory4a[307 ] = 3'd2;
    assign memory4a[308 ] = 3'd2;
    assign memory4a[309 ] = 3'd1;
    assign memory4a[310 ] = 3'd0;
    assign memory4a[311 ] = 3'd1;
    assign memory4a[312 ] = 3'd2;
    assign memory4a[313 ] = 3'd2;
    assign memory4a[314 ] = 3'd2;
    assign memory4a[315 ] = 3'd2;
    assign memory4a[316 ] = 3'd2;
    assign memory4a[317 ] = 3'd2;
    assign memory4a[318 ] = 3'd2;
    assign memory4a[319 ] = 3'd2;
    assign memory4a[320 ] = 3'd2;
    assign memory4a[321 ] = 3'd4;
    assign memory4a[322 ] = 3'd5;
    assign memory4a[323 ] = 3'd5;
    assign memory4a[324 ] = 3'd5;
    assign memory4a[325 ] = 3'd5;
    assign memory4a[326 ] = 3'd4;
    assign memory4a[327 ] = 3'd2;
    assign memory4a[328 ] = 3'd2;
    assign memory4a[329 ] = 3'd1;
    assign memory4a[330 ] = 3'd0;
    assign memory4a[331 ] = 3'd1;
    assign memory4a[332 ] = 3'd2;
    assign memory4a[333 ] = 3'd2;
    assign memory4a[334 ] = 3'd2;
    assign memory4a[335 ] = 3'd2;
    assign memory4a[336 ] = 3'd2;
    assign memory4a[337 ] = 3'd2;
    assign memory4a[338 ] = 3'd2;
    assign memory4a[339 ] = 3'd2;
    assign memory4a[340 ] = 3'd1;
    assign memory4a[341 ] = 3'd0;
    assign memory4a[342 ] = 3'd1;
    assign memory4a[343 ] = 3'd2;
    assign memory4a[344 ] = 3'd2;
    assign memory4a[345 ] = 3'd2;
    assign memory4a[346 ] = 3'd2;
    assign memory4a[347 ] = 3'd2;
    assign memory4a[348 ] = 3'd2;
    assign memory4a[349 ] = 3'd2;
    assign memory4a[350 ] = 3'd2;
    assign memory4a[351 ] = 3'd2;
    assign memory4a[352 ] = 3'd2;
    assign memory4a[353 ] = 3'd4;
    assign memory4a[354 ] = 3'd5;
    assign memory4a[355 ] = 3'd5;
    assign memory4a[356 ] = 3'd5;
    assign memory4a[357 ] = 3'd5;
    assign memory4a[358 ] = 3'd4;
    assign memory4a[359 ] = 3'd2;
    assign memory4a[360 ] = 3'd2;
    assign memory4a[361 ] = 3'd2;
    assign memory4a[362 ] = 3'd1;
    assign memory4a[363 ] = 3'd0;
    assign memory4a[364 ] = 3'd1;
    assign memory4a[365 ] = 3'd2;
    assign memory4a[366 ] = 3'd2;
    assign memory4a[367 ] = 3'd2;
    assign memory4a[368 ] = 3'd2;
    assign memory4a[369 ] = 3'd2;
    assign memory4a[370 ] = 3'd2;
    assign memory4a[371 ] = 3'd1;
    assign memory4a[372 ] = 3'd0;
    assign memory4a[373 ] = 3'd1;
    assign memory4a[374 ] = 3'd2;
    assign memory4a[375 ] = 3'd2;
    assign memory4a[376 ] = 3'd2;
    assign memory4a[377 ] = 3'd2;
    assign memory4a[378 ] = 3'd2;
    assign memory4a[379 ] = 3'd2;
    assign memory4a[380 ] = 3'd2;
    assign memory4a[381 ] = 3'd2;
    assign memory4a[382 ] = 3'd2;
    assign memory4a[383 ] = 3'd2;
    assign memory4a[384 ] = 3'd2;
    assign memory4a[385 ] = 3'd4;
    assign memory4a[386 ] = 3'd4;
    assign memory4a[387 ] = 3'd4;
    assign memory4a[388 ] = 3'd4;
    assign memory4a[389 ] = 3'd4;
    assign memory4a[390 ] = 3'd4;
    assign memory4a[391 ] = 3'd2;
    assign memory4a[392 ] = 3'd2;
    assign memory4a[393 ] = 3'd2;
    assign memory4a[394 ] = 3'd2;
    assign memory4a[395 ] = 3'd1;
    assign memory4a[396 ] = 3'd0;
    assign memory4a[397 ] = 3'd1;
    assign memory4a[398 ] = 3'd2;
    assign memory4a[399 ] = 3'd2;
    assign memory4a[400 ] = 3'd2;
    assign memory4a[401 ] = 3'd2;
    assign memory4a[402 ] = 3'd1;
    assign memory4a[403 ] = 3'd0;
    assign memory4a[404 ] = 3'd1;
    assign memory4a[405 ] = 3'd2;
    assign memory4a[406 ] = 3'd2;
    assign memory4a[407 ] = 3'd2;
    assign memory4a[408 ] = 3'd2;
    assign memory4a[409 ] = 3'd2;
    assign memory4a[410 ] = 3'd2;
    assign memory4a[411 ] = 3'd2;
    assign memory4a[412 ] = 3'd2;
    assign memory4a[413 ] = 3'd2;
    assign memory4a[414 ] = 3'd2;
    assign memory4a[415 ] = 3'd2;
    assign memory4a[416 ] = 3'd2;
    assign memory4a[417 ] = 3'd2;
    assign memory4a[418 ] = 3'd2;
    assign memory4a[419 ] = 3'd2;
    assign memory4a[420 ] = 3'd2;
    assign memory4a[421 ] = 3'd2;
    assign memory4a[422 ] = 3'd2;
    assign memory4a[423 ] = 3'd2;
    assign memory4a[424 ] = 3'd2;
    assign memory4a[425 ] = 3'd2;
    assign memory4a[426 ] = 3'd2;
    assign memory4a[427 ] = 3'd2;
    assign memory4a[428 ] = 3'd1;
    assign memory4a[429 ] = 3'd0;
    assign memory4a[430 ] = 3'd1;
    assign memory4a[431 ] = 3'd2;
    assign memory4a[432 ] = 3'd2;
    assign memory4a[433 ] = 3'd1;
    assign memory4a[434 ] = 3'd0;
    assign memory4a[435 ] = 3'd1;
    assign memory4a[436 ] = 3'd2;
    assign memory4a[437 ] = 3'd2;
    assign memory4a[438 ] = 3'd2;
    assign memory4a[439 ] = 3'd2;
    assign memory4a[440 ] = 3'd2;
    assign memory4a[441 ] = 3'd2;
    assign memory4a[442 ] = 3'd2;
    assign memory4a[443 ] = 3'd2;
    assign memory4a[444 ] = 3'd2;
    assign memory4a[445 ] = 3'd2;
    assign memory4a[446 ] = 3'd2;
    assign memory4a[447 ] = 3'd2;
    assign memory4a[448 ] = 3'd2;
    assign memory4a[449 ] = 3'd2;
    assign memory4a[450 ] = 3'd2;
    assign memory4a[451 ] = 3'd2;
    assign memory4a[452 ] = 3'd2;
    assign memory4a[453 ] = 3'd2;
    assign memory4a[454 ] = 3'd2;
    assign memory4a[455 ] = 3'd2;
    assign memory4a[456 ] = 3'd2;
    assign memory4a[457 ] = 3'd2;
    assign memory4a[458 ] = 3'd2;
    assign memory4a[459 ] = 3'd2;
    assign memory4a[460 ] = 3'd2;
    assign memory4a[461 ] = 3'd1;
    assign memory4a[462 ] = 3'd0;
    assign memory4a[463 ] = 3'd1;
    assign memory4a[464 ] = 3'd1;
    assign memory4a[465 ] = 3'd0;
    assign memory4a[466 ] = 3'd1;
    assign memory4a[467 ] = 3'd2;
    assign memory4a[468 ] = 3'd2;
    assign memory4a[469 ] = 3'd2;
    assign memory4a[470 ] = 3'd2;
    assign memory4a[471 ] = 3'd2;
    assign memory4a[472 ] = 3'd2;
    assign memory4a[473 ] = 3'd2;
    assign memory4a[474 ] = 3'd2;
    assign memory4a[475 ] = 3'd2;
    assign memory4a[476 ] = 3'd2;
    assign memory4a[477 ] = 3'd2;
    assign memory4a[478 ] = 3'd2;
    assign memory4a[479 ] = 3'd2;
    assign memory4a[480 ] = 3'd2;
    assign memory4a[481 ] = 3'd2;
    assign memory4a[482 ] = 3'd2;
    assign memory4a[483 ] = 3'd2;
    assign memory4a[484 ] = 3'd2;
    assign memory4a[485 ] = 3'd2;
    assign memory4a[486 ] = 3'd2;
    assign memory4a[487 ] = 3'd2;
    assign memory4a[488 ] = 3'd2;
    assign memory4a[489 ] = 3'd2;
    assign memory4a[490 ] = 3'd2;
    assign memory4a[491 ] = 3'd2;
    assign memory4a[492 ] = 3'd2;
    assign memory4a[493 ] = 3'd2;
    assign memory4a[494 ] = 3'd1;
    assign memory4a[495 ] = 3'd0;
    assign memory4a[496 ] = 3'd0;
    assign memory4a[497 ] = 3'd1;
    assign memory4a[498 ] = 3'd2;
    assign memory4a[499 ] = 3'd2;
    assign memory4a[500 ] = 3'd2;
    assign memory4a[501 ] = 3'd2;
    assign memory4a[502 ] = 3'd2;
    assign memory4a[503 ] = 3'd2;
    assign memory4a[504 ] = 3'd2;
    assign memory4a[505 ] = 3'd2;
    assign memory4a[506 ] = 3'd2;
    assign memory4a[507 ] = 3'd2;
    assign memory4a[508 ] = 3'd2;
    assign memory4a[509 ] = 3'd2;
    assign memory4a[510 ] = 3'd2;
    assign memory4a[511 ] = 3'd2;
    assign memory4a[512 ] = 3'd2;
    assign memory4a[513 ] = 3'd2;
    assign memory4a[514 ] = 3'd2;
    assign memory4a[515 ] = 3'd2;
    assign memory4a[516 ] = 3'd2;
    assign memory4a[517 ] = 3'd2;
    assign memory4a[518 ] = 3'd2;
    assign memory4a[519 ] = 3'd2;
    assign memory4a[520 ] = 3'd2;
    assign memory4a[521 ] = 3'd2;
    assign memory4a[522 ] = 3'd2;
    assign memory4a[523 ] = 3'd2;
    assign memory4a[524 ] = 3'd2;
    assign memory4a[525 ] = 3'd2;
    assign memory4a[526 ] = 3'd1;
    assign memory4a[527 ] = 3'd0;
    assign memory4a[528 ] = 3'd0;
    assign memory4a[529 ] = 3'd1;
    assign memory4a[530 ] = 3'd2;
    assign memory4a[531 ] = 3'd2;
    assign memory4a[532 ] = 3'd2;
    assign memory4a[533 ] = 3'd2;
    assign memory4a[534 ] = 3'd2;
    assign memory4a[535 ] = 3'd2;
    assign memory4a[536 ] = 3'd2;
    assign memory4a[537 ] = 3'd2;
    assign memory4a[538 ] = 3'd2;
    assign memory4a[539 ] = 3'd2;
    assign memory4a[540 ] = 3'd2;
    assign memory4a[541 ] = 3'd2;
    assign memory4a[542 ] = 3'd2;
    assign memory4a[543 ] = 3'd2;
    assign memory4a[544 ] = 3'd2;
    assign memory4a[545 ] = 3'd2;
    assign memory4a[546 ] = 3'd2;
    assign memory4a[547 ] = 3'd2;
    assign memory4a[548 ] = 3'd2;
    assign memory4a[549 ] = 3'd2;
    assign memory4a[550 ] = 3'd2;
    assign memory4a[551 ] = 3'd2;
    assign memory4a[552 ] = 3'd2;
    assign memory4a[553 ] = 3'd2;
    assign memory4a[554 ] = 3'd2;
    assign memory4a[555 ] = 3'd2;
    assign memory4a[556 ] = 3'd2;
    assign memory4a[557 ] = 3'd1;
    assign memory4a[558 ] = 3'd0;
    assign memory4a[559 ] = 3'd1;
    assign memory4a[560 ] = 3'd1;
    assign memory4a[561 ] = 3'd0;
    assign memory4a[562 ] = 3'd1;
    assign memory4a[563 ] = 3'd2;
    assign memory4a[564 ] = 3'd2;
    assign memory4a[565 ] = 3'd2;
    assign memory4a[566 ] = 3'd2;
    assign memory4a[567 ] = 3'd2;
    assign memory4a[568 ] = 3'd2;
    assign memory4a[569 ] = 3'd2;
    assign memory4a[570 ] = 3'd2;
    assign memory4a[571 ] = 3'd2;
    assign memory4a[572 ] = 3'd2;
    assign memory4a[573 ] = 3'd2;
    assign memory4a[574 ] = 3'd2;
    assign memory4a[575 ] = 3'd2;
    assign memory4a[576 ] = 3'd2;
    assign memory4a[577 ] = 3'd2;
    assign memory4a[578 ] = 3'd2;
    assign memory4a[579 ] = 3'd2;
    assign memory4a[580 ] = 3'd2;
    assign memory4a[581 ] = 3'd2;
    assign memory4a[582 ] = 3'd2;
    assign memory4a[583 ] = 3'd2;
    assign memory4a[584 ] = 3'd2;
    assign memory4a[585 ] = 3'd2;
    assign memory4a[586 ] = 3'd2;
    assign memory4a[587 ] = 3'd2;
    assign memory4a[588 ] = 3'd1;
    assign memory4a[589 ] = 3'd0;
    assign memory4a[590 ] = 3'd1;
    assign memory4a[591 ] = 3'd2;
    assign memory4a[592 ] = 3'd2;
    assign memory4a[593 ] = 3'd1;
    assign memory4a[594 ] = 3'd0;
    assign memory4a[595 ] = 3'd1;
    assign memory4a[596 ] = 3'd2;
    assign memory4a[597 ] = 3'd2;
    assign memory4a[598 ] = 3'd2;
    assign memory4a[599 ] = 3'd2;
    assign memory4a[600 ] = 3'd2;
    assign memory4a[601 ] = 3'd2;
    assign memory4a[602 ] = 3'd2;
    assign memory4a[603 ] = 3'd2;
    assign memory4a[604 ] = 3'd2;
    assign memory4a[605 ] = 3'd2;
    assign memory4a[606 ] = 3'd2;
    assign memory4a[607 ] = 3'd2;
    assign memory4a[608 ] = 3'd2;
    assign memory4a[609 ] = 3'd2;
    assign memory4a[610 ] = 3'd2;
    assign memory4a[611 ] = 3'd2;
    assign memory4a[612 ] = 3'd2;
    assign memory4a[613 ] = 3'd2;
    assign memory4a[614 ] = 3'd2;
    assign memory4a[615 ] = 3'd2;
    assign memory4a[616 ] = 3'd2;
    assign memory4a[617 ] = 3'd2;
    assign memory4a[618 ] = 3'd2;
    assign memory4a[619 ] = 3'd1;
    assign memory4a[620 ] = 3'd0;
    assign memory4a[621 ] = 3'd1;
    assign memory4a[622 ] = 3'd2;
    assign memory4a[623 ] = 3'd2;
    assign memory4a[624 ] = 3'd2;
    assign memory4a[625 ] = 3'd2;
    assign memory4a[626 ] = 3'd1;
    assign memory4a[627 ] = 3'd0;
    assign memory4a[628 ] = 3'd1;
    assign memory4a[629 ] = 3'd2;
    assign memory4a[630 ] = 3'd2;
    assign memory4a[631 ] = 3'd2;
    assign memory4a[632 ] = 3'd2;
    assign memory4a[633 ] = 3'd2;
    assign memory4a[634 ] = 3'd2;
    assign memory4a[635 ] = 3'd2;
    assign memory4a[636 ] = 3'd2;
    assign memory4a[637 ] = 3'd2;
    assign memory4a[638 ] = 3'd2;
    assign memory4a[639 ] = 3'd2;
    assign memory4a[640 ] = 3'd2;
    assign memory4a[641 ] = 3'd2;
    assign memory4a[642 ] = 3'd2;
    assign memory4a[643 ] = 3'd2;
    assign memory4a[644 ] = 3'd2;
    assign memory4a[645 ] = 3'd2;
    assign memory4a[646 ] = 3'd2;
    assign memory4a[647 ] = 3'd2;
    assign memory4a[648 ] = 3'd2;
    assign memory4a[649 ] = 3'd2;
    assign memory4a[650 ] = 3'd1;
    assign memory4a[651 ] = 3'd0;
    assign memory4a[652 ] = 3'd1;
    assign memory4a[653 ] = 3'd2;
    assign memory4a[654 ] = 3'd2;
    assign memory4a[655 ] = 3'd2;
    assign memory4a[656 ] = 3'd2;
    assign memory4a[657 ] = 3'd2;
    assign memory4a[658 ] = 3'd2;
    assign memory4a[659 ] = 3'd1;
    assign memory4a[660 ] = 3'd0;
    assign memory4a[661 ] = 3'd1;
    assign memory4a[662 ] = 3'd2;
    assign memory4a[663 ] = 3'd2;
    assign memory4a[664 ] = 3'd2;
    assign memory4a[665 ] = 3'd2;
    assign memory4a[666 ] = 3'd2;
    assign memory4a[667 ] = 3'd2;
    assign memory4a[668 ] = 3'd2;
    assign memory4a[669 ] = 3'd2;
    assign memory4a[670 ] = 3'd2;
    assign memory4a[671 ] = 3'd2;
    assign memory4a[672 ] = 3'd2;
    assign memory4a[673 ] = 3'd2;
    assign memory4a[674 ] = 3'd2;
    assign memory4a[675 ] = 3'd2;
    assign memory4a[676 ] = 3'd2;
    assign memory4a[677 ] = 3'd2;
    assign memory4a[678 ] = 3'd2;
    assign memory4a[679 ] = 3'd2;
    assign memory4a[680 ] = 3'd2;
    assign memory4a[681 ] = 3'd1;
    assign memory4a[682 ] = 3'd0;
    assign memory4a[683 ] = 3'd1;
    assign memory4a[684 ] = 3'd2;
    assign memory4a[685 ] = 3'd2;
    assign memory4a[686 ] = 3'd2;
    assign memory4a[687 ] = 3'd2;
    assign memory4a[688 ] = 3'd2;
    assign memory4a[689 ] = 3'd2;
    assign memory4a[690 ] = 3'd2;
    assign memory4a[691 ] = 3'd2;
    assign memory4a[692 ] = 3'd1;
    assign memory4a[693 ] = 3'd0;
    assign memory4a[694 ] = 3'd2;
    assign memory4a[695 ] = 3'd2;
    assign memory4a[696 ] = 3'd2;
    assign memory4a[697 ] = 3'd2;
    assign memory4a[698 ] = 3'd2;
    assign memory4a[699 ] = 3'd2;
    assign memory4a[700 ] = 3'd2;
    assign memory4a[701 ] = 3'd2;
    assign memory4a[702 ] = 3'd2;
    assign memory4a[703 ] = 3'd2;
    assign memory4a[704 ] = 3'd2;
    assign memory4a[705 ] = 3'd2;
    assign memory4a[706 ] = 3'd2;
    assign memory4a[707 ] = 3'd2;
    assign memory4a[708 ] = 3'd2;
    assign memory4a[709 ] = 3'd2;
    assign memory4a[710 ] = 3'd2;
    assign memory4a[711 ] = 3'd2;
    assign memory4a[712 ] = 3'd1;
    assign memory4a[713 ] = 3'd0;
    assign memory4a[714 ] = 3'd1;
    assign memory4a[715 ] = 3'd2;
    assign memory4a[716 ] = 3'd2;
    assign memory4a[717 ] = 3'd2;
    assign memory4a[718 ] = 3'd2;
    assign memory4a[719 ] = 3'd2;
    assign memory4a[720 ] = 3'd2;
    assign memory4a[721 ] = 3'd2;
    assign memory4a[722 ] = 3'd2;
    assign memory4a[723 ] = 3'd2;
    assign memory4a[724 ] = 3'd2;
    assign memory4a[725 ] = 3'd1;
    assign memory4a[726 ] = 3'd0;
    assign memory4a[727 ] = 3'd1;
    assign memory4a[728 ] = 3'd2;
    assign memory4a[729 ] = 3'd2;
    assign memory4a[730 ] = 3'd2;
    assign memory4a[731 ] = 3'd2;
    assign memory4a[732 ] = 3'd2;
    assign memory4a[733 ] = 3'd2;
    assign memory4a[734 ] = 3'd2;
    assign memory4a[735 ] = 3'd2;
    assign memory4a[736 ] = 3'd2;
    assign memory4a[737 ] = 3'd2;
    assign memory4a[738 ] = 3'd2;
    assign memory4a[739 ] = 3'd2;
    assign memory4a[740 ] = 3'd2;
    assign memory4a[741 ] = 3'd2;
    assign memory4a[742 ] = 3'd2;
    assign memory4a[743 ] = 3'd1;
    assign memory4a[744 ] = 3'd0;
    assign memory4a[745 ] = 3'd1;
    assign memory4a[746 ] = 3'd2;
    assign memory4a[747 ] = 3'd2;
    assign memory4a[748 ] = 3'd2;
    assign memory4a[749 ] = 3'd2;
    assign memory4a[750 ] = 3'd2;
    assign memory4a[751 ] = 3'd2;
    assign memory4a[752 ] = 3'd2;
    assign memory4a[753 ] = 3'd2;
    assign memory4a[754 ] = 3'd2;
    assign memory4a[755 ] = 3'd2;
    assign memory4a[756 ] = 3'd2;
    assign memory4a[757 ] = 3'd2;
    assign memory4a[758 ] = 3'd1;
    assign memory4a[759 ] = 3'd0;
    assign memory4a[760 ] = 3'd1;
    assign memory4a[761 ] = 3'd2;
    assign memory4a[762 ] = 3'd2;
    assign memory4a[763 ] = 3'd2;
    assign memory4a[764 ] = 3'd2;
    assign memory4a[765 ] = 3'd2;
    assign memory4a[766 ] = 3'd2;
    assign memory4a[767 ] = 3'd2;
    assign memory4a[768 ] = 3'd2;
    assign memory4a[769 ] = 3'd2;
    assign memory4a[770 ] = 3'd2;
    assign memory4a[771 ] = 3'd2;
    assign memory4a[772 ] = 3'd2;
    assign memory4a[773 ] = 3'd2;
    assign memory4a[774 ] = 3'd1;
    assign memory4a[775 ] = 3'd0;
    assign memory4a[776 ] = 3'd1;
    assign memory4a[777 ] = 3'd2;
    assign memory4a[778 ] = 3'd2;
    assign memory4a[779 ] = 3'd2;
    assign memory4a[780 ] = 3'd2;
    assign memory4a[781 ] = 3'd2;
    assign memory4a[782 ] = 3'd2;
    assign memory4a[783 ] = 3'd2;
    assign memory4a[784 ] = 3'd2;
    assign memory4a[785 ] = 3'd2;
    assign memory4a[786 ] = 3'd2;
    assign memory4a[787 ] = 3'd2;
    assign memory4a[788 ] = 3'd2;
    assign memory4a[789 ] = 3'd2;
    assign memory4a[790 ] = 3'd2;
    assign memory4a[791 ] = 3'd1;
    assign memory4a[792 ] = 3'd0;
    assign memory4a[793 ] = 3'd3;
    assign memory4a[794 ] = 3'd2;
    assign memory4a[795 ] = 3'd2;
    assign memory4a[796 ] = 3'd2;
    assign memory4a[797 ] = 3'd2;
    assign memory4a[798 ] = 3'd2;
    assign memory4a[799 ] = 3'd2;
    assign memory4a[800 ] = 3'd2;
    assign memory4a[801 ] = 3'd2;
    assign memory4a[802 ] = 3'd2;
    assign memory4a[803 ] = 3'd2;
    assign memory4a[804 ] = 3'd2;
    assign memory4a[805 ] = 3'd1;
    assign memory4a[806 ] = 3'd0;
    assign memory4a[807 ] = 3'd1;
    assign memory4a[808 ] = 3'd2;
    assign memory4a[809 ] = 3'd2;
    assign memory4a[810 ] = 3'd2;
    assign memory4a[811 ] = 3'd2;
    assign memory4a[812 ] = 3'd2;
    assign memory4a[813 ] = 3'd2;
    assign memory4a[814 ] = 3'd2;
    assign memory4a[815 ] = 3'd2;
    assign memory4a[816 ] = 3'd2;
    assign memory4a[817 ] = 3'd2;
    assign memory4a[818 ] = 3'd2;
    assign memory4a[819 ] = 3'd2;
    assign memory4a[820 ] = 3'd2;
    assign memory4a[821 ] = 3'd2;
    assign memory4a[822 ] = 3'd4;
    assign memory4a[823 ] = 3'd2;
    assign memory4a[824 ] = 3'd3;
    assign memory4a[825 ] = 3'd3;
    assign memory4a[826 ] = 3'd2;
    assign memory4a[827 ] = 3'd4;
    assign memory4a[828 ] = 3'd2;
    assign memory4a[829 ] = 3'd2;
    assign memory4a[830 ] = 3'd2;
    assign memory4a[831 ] = 3'd2;
    assign memory4a[832 ] = 3'd2;
    assign memory4a[833 ] = 3'd2;
    assign memory4a[834 ] = 3'd2;
    assign memory4a[835 ] = 3'd2;
    assign memory4a[836 ] = 3'd1;
    assign memory4a[837 ] = 3'd0;
    assign memory4a[838 ] = 3'd1;
    assign memory4a[839 ] = 3'd2;
    assign memory4a[840 ] = 3'd2;
    assign memory4a[841 ] = 3'd2;
    assign memory4a[842 ] = 3'd2;
    assign memory4a[843 ] = 3'd2;
    assign memory4a[844 ] = 3'd2;
    assign memory4a[845 ] = 3'd2;
    assign memory4a[846 ] = 3'd2;
    assign memory4a[847 ] = 3'd2;
    assign memory4a[848 ] = 3'd2;
    assign memory4a[849 ] = 3'd2;
    assign memory4a[850 ] = 3'd2;
    assign memory4a[851 ] = 3'd2;
    assign memory4a[852 ] = 3'd2;
    assign memory4a[853 ] = 3'd2;
    assign memory4a[854 ] = 3'd4;
    assign memory4a[855 ] = 3'd2;
    assign memory4a[856 ] = 3'd3;
    assign memory4a[857 ] = 3'd3;
    assign memory4a[858 ] = 3'd0;
    assign memory4a[859 ] = 3'd4;
    assign memory4a[860 ] = 3'd2;
    assign memory4a[861 ] = 3'd2;
    assign memory4a[862 ] = 3'd2;
    assign memory4a[863 ] = 3'd2;
    assign memory4a[864 ] = 3'd2;
    assign memory4a[865 ] = 3'd2;
    assign memory4a[866 ] = 3'd2;
    assign memory4a[867 ] = 3'd1;
    assign memory4a[868 ] = 3'd0;
    assign memory4a[869 ] = 3'd1;
    assign memory4a[870 ] = 3'd2;
    assign memory4a[871 ] = 3'd2;
    assign memory4a[872 ] = 3'd2;
    assign memory4a[873 ] = 3'd2;
    assign memory4a[874 ] = 3'd2;
    assign memory4a[875 ] = 3'd2;
    assign memory4a[876 ] = 3'd2;
    assign memory4a[877 ] = 3'd2;
    assign memory4a[878 ] = 3'd2;
    assign memory4a[879 ] = 3'd2;
    assign memory4a[880 ] = 3'd2;
    assign memory4a[881 ] = 3'd2;
    assign memory4a[882 ] = 3'd2;
    assign memory4a[883 ] = 3'd2;
    assign memory4a[884 ] = 3'd2;
    assign memory4a[885 ] = 3'd2;
    assign memory4a[886 ] = 3'd4;
    assign memory4a[887 ] = 3'd5;
    assign memory4a[888 ] = 3'd5;
    assign memory4a[889 ] = 3'd5;
    assign memory4a[890 ] = 3'd5;
    assign memory4a[891 ] = 3'd4;
    assign memory4a[892 ] = 3'd1;
    assign memory4a[893 ] = 3'd2;
    assign memory4a[894 ] = 3'd2;
    assign memory4a[895 ] = 3'd2;
    assign memory4a[896 ] = 3'd2;
    assign memory4a[897 ] = 3'd2;
    assign memory4a[898 ] = 3'd1;
    assign memory4a[899 ] = 3'd0;
    assign memory4a[900 ] = 3'd1;
    assign memory4a[901 ] = 3'd2;
    assign memory4a[902 ] = 3'd2;
    assign memory4a[903 ] = 3'd2;
    assign memory4a[904 ] = 3'd2;
    assign memory4a[905 ] = 3'd2;
    assign memory4a[906 ] = 3'd2;
    assign memory4a[907 ] = 3'd2;
    assign memory4a[908 ] = 3'd2;
    assign memory4a[909 ] = 3'd2;
    assign memory4a[910 ] = 3'd2;
    assign memory4a[911 ] = 3'd2;
    assign memory4a[912 ] = 3'd2;
    assign memory4a[913 ] = 3'd2;
    assign memory4a[914 ] = 3'd2;
    assign memory4a[915 ] = 3'd2;
    assign memory4a[916 ] = 3'd2;
    assign memory4a[917 ] = 3'd2;
    assign memory4a[918 ] = 3'd4;
    assign memory4a[919 ] = 3'd5;
    assign memory4a[920 ] = 3'd5;
    assign memory4a[921 ] = 3'd5;
    assign memory4a[922 ] = 3'd5;
    assign memory4a[923 ] = 3'd4;
    assign memory4a[924 ] = 3'd0;
    assign memory4a[925 ] = 3'd1;
    assign memory4a[926 ] = 3'd2;
    assign memory4a[927 ] = 3'd2;
    assign memory4a[928 ] = 3'd2;
    assign memory4a[929 ] = 3'd1;
    assign memory4a[930 ] = 3'd0;
    assign memory4a[931 ] = 3'd1;
    assign memory4a[932 ] = 3'd2;
    assign memory4a[933 ] = 3'd2;
    assign memory4a[934 ] = 3'd2;
    assign memory4a[935 ] = 3'd2;
    assign memory4a[936 ] = 3'd2;
    assign memory4a[937 ] = 3'd2;
    assign memory4a[938 ] = 3'd2;
    assign memory4a[939 ] = 3'd2;
    assign memory4a[940 ] = 3'd2;
    assign memory4a[941 ] = 3'd2;
    assign memory4a[942 ] = 3'd2;
    assign memory4a[943 ] = 3'd2;
    assign memory4a[944 ] = 3'd2;
    assign memory4a[945 ] = 3'd2;
    assign memory4a[946 ] = 3'd2;
    assign memory4a[947 ] = 3'd2;
    assign memory4a[948 ] = 3'd2;
    assign memory4a[949 ] = 3'd2;
    assign memory4a[950 ] = 3'd4;
    assign memory4a[951 ] = 3'd5;
    assign memory4a[952 ] = 3'd5;
    assign memory4a[953 ] = 3'd5;
    assign memory4a[954 ] = 3'd5;
    assign memory4a[955 ] = 3'd4;
    assign memory4a[956 ] = 3'd1;
    assign memory4a[957 ] = 3'd0;
    assign memory4a[958 ] = 3'd1;
    assign memory4a[959 ] = 3'd2;
    assign memory4a[960 ] = 3'd1;
    assign memory4a[961 ] = 3'd0;
    assign memory4a[962 ] = 3'd1;
    assign memory4a[963 ] = 3'd2;
    assign memory4a[964 ] = 3'd2;
    assign memory4a[965 ] = 3'd2;
    assign memory4a[966 ] = 3'd2;
    assign memory4a[967 ] = 3'd2;
    assign memory4a[968 ] = 3'd2;
    assign memory4a[969 ] = 3'd2;
    assign memory4a[970 ] = 3'd2;
    assign memory4a[971 ] = 3'd2;
    assign memory4a[972 ] = 3'd2;
    assign memory4a[973 ] = 3'd2;
    assign memory4a[974 ] = 3'd2;
    assign memory4a[975 ] = 3'd2;
    assign memory4a[976 ] = 3'd2;
    assign memory4a[977 ] = 3'd2;
    assign memory4a[978 ] = 3'd2;
    assign memory4a[979 ] = 3'd2;
    assign memory4a[980 ] = 3'd2;
    assign memory4a[981 ] = 3'd2;
    assign memory4a[982 ] = 3'd4;
    assign memory4a[983 ] = 3'd5;
    assign memory4a[984 ] = 3'd5;
    assign memory4a[985 ] = 3'd5;
    assign memory4a[986 ] = 3'd5;
    assign memory4a[987 ] = 3'd4;
    assign memory4a[988 ] = 3'd2;
    assign memory4a[989 ] = 3'd1;
    assign memory4a[990 ] = 3'd0;
    assign memory4a[991 ] = 3'd1;
    assign memory4a[992 ] = 3'd0;
    assign memory4a[993 ] = 3'd1;
    assign memory4a[994 ] = 3'd2;
    assign memory4a[995 ] = 3'd2;
    assign memory4a[996 ] = 3'd2;
    assign memory4a[997 ] = 3'd2;
    assign memory4a[998 ] = 3'd2;
    assign memory4a[999 ] = 3'd2;
    assign memory4a[1000] = 3'd2;
    assign memory4a[1001] = 3'd2;
    assign memory4a[1002] = 3'd2;
    assign memory4a[1003] = 3'd2;
    assign memory4a[1004] = 3'd2;
    assign memory4a[1005] = 3'd2;
    assign memory4a[1006] = 3'd2;
    assign memory4a[1007] = 3'd2;
    assign memory4a[1008] = 3'd2;
    assign memory4a[1009] = 3'd2;
    assign memory4a[1010] = 3'd2;
    assign memory4a[1011] = 3'd2;
    assign memory4a[1012] = 3'd2;
    assign memory4a[1013] = 3'd2;
    assign memory4a[1014] = 3'd4;
    assign memory4a[1015] = 3'd4;
    assign memory4a[1016] = 3'd4;
    assign memory4a[1017] = 3'd4;
    assign memory4a[1018] = 3'd4;
    assign memory4a[1019] = 3'd4;
    assign memory4a[1020] = 3'd2;
    assign memory4a[1021] = 3'd2;
    assign memory4a[1022] = 3'd1;
    assign memory4a[1023] = 3'd0;

    assign memory4b[0   ] = 3'd0;
    assign memory4b[1   ] = 3'd0;
    assign memory4b[2   ] = 3'd0;
    assign memory4b[3   ] = 3'd0;
    assign memory4b[4   ] = 3'd0;
    assign memory4b[5   ] = 3'd0;
    assign memory4b[6   ] = 3'd0;
    assign memory4b[7   ] = 3'd0;
    assign memory4b[8   ] = 3'd0;
    assign memory4b[9   ] = 3'd0;
    assign memory4b[10  ] = 3'd0;
    assign memory4b[11  ] = 3'd0;
    assign memory4b[12  ] = 3'd0;
    assign memory4b[13  ] = 3'd0;
    assign memory4b[14  ] = 3'd0;
    assign memory4b[15  ] = 3'd0;
    assign memory4b[16  ] = 3'd0;
    assign memory4b[17  ] = 3'd0;
    assign memory4b[18  ] = 3'd0;
    assign memory4b[19  ] = 3'd0;
    assign memory4b[20  ] = 3'd0;
    assign memory4b[21  ] = 3'd0;
    assign memory4b[22  ] = 3'd0;
    assign memory4b[23  ] = 3'd0;
    assign memory4b[24  ] = 3'd0;
    assign memory4b[25  ] = 3'd0;
    assign memory4b[26  ] = 3'd0;
    assign memory4b[27  ] = 3'd0;
    assign memory4b[28  ] = 3'd0;
    assign memory4b[29  ] = 3'd0;
    assign memory4b[30  ] = 3'd0;
    assign memory4b[31  ] = 3'd0;
    assign memory4b[32  ] = 3'd0;
    assign memory4b[33  ] = 3'd1;
    assign memory4b[34  ] = 3'd1;
    assign memory4b[35  ] = 3'd1;
    assign memory4b[36  ] = 3'd1;
    assign memory4b[37  ] = 3'd1;
    assign memory4b[38  ] = 3'd1;
    assign memory4b[39  ] = 3'd1;
    assign memory4b[40  ] = 3'd1;
    assign memory4b[41  ] = 3'd1;
    assign memory4b[42  ] = 3'd1;
    assign memory4b[43  ] = 3'd1;
    assign memory4b[44  ] = 3'd1;
    assign memory4b[45  ] = 3'd1;
    assign memory4b[46  ] = 3'd1;
    assign memory4b[47  ] = 3'd1;
    assign memory4b[48  ] = 3'd1;
    assign memory4b[49  ] = 3'd1;
    assign memory4b[50  ] = 3'd1;
    assign memory4b[51  ] = 3'd1;
    assign memory4b[52  ] = 3'd1;
    assign memory4b[53  ] = 3'd1;
    assign memory4b[54  ] = 3'd1;
    assign memory4b[55  ] = 3'd1;
    assign memory4b[56  ] = 3'd1;
    assign memory4b[57  ] = 3'd1;
    assign memory4b[58  ] = 3'd1;
    assign memory4b[59  ] = 3'd1;
    assign memory4b[60  ] = 3'd1;
    assign memory4b[61  ] = 3'd1;
    assign memory4b[62  ] = 3'd1;
    assign memory4b[63  ] = 3'd0;
    assign memory4b[64  ] = 3'd0;
    assign memory4b[65  ] = 3'd1;
    assign memory4b[66  ] = 3'd1;
    assign memory4b[67  ] = 3'd1;
    assign memory4b[68  ] = 3'd1;
    assign memory4b[69  ] = 3'd1;
    assign memory4b[70  ] = 3'd1;
    assign memory4b[71  ] = 3'd1;
    assign memory4b[72  ] = 3'd1;
    assign memory4b[73  ] = 3'd1;
    assign memory4b[74  ] = 3'd1;
    assign memory4b[75  ] = 3'd1;
    assign memory4b[76  ] = 3'd1;
    assign memory4b[77  ] = 3'd1;
    assign memory4b[78  ] = 3'd1;
    assign memory4b[79  ] = 3'd1;
    assign memory4b[80  ] = 3'd1;
    assign memory4b[81  ] = 3'd1;
    assign memory4b[82  ] = 3'd1;
    assign memory4b[83  ] = 3'd1;
    assign memory4b[84  ] = 3'd1;
    assign memory4b[85  ] = 3'd1;
    assign memory4b[86  ] = 3'd1;
    assign memory4b[87  ] = 3'd1;
    assign memory4b[88  ] = 3'd1;
    assign memory4b[89  ] = 3'd1;
    assign memory4b[90  ] = 3'd1;
    assign memory4b[91  ] = 3'd1;
    assign memory4b[92  ] = 3'd1;
    assign memory4b[93  ] = 3'd1;
    assign memory4b[94  ] = 3'd1;
    assign memory4b[95  ] = 3'd0;
    assign memory4b[96  ] = 3'd0;
    assign memory4b[97  ] = 3'd1;
    assign memory4b[98  ] = 3'd1;
    assign memory4b[99  ] = 3'd2;
    assign memory4b[100 ] = 3'd2;
    assign memory4b[101 ] = 3'd2;
    assign memory4b[102 ] = 3'd1;
    assign memory4b[103 ] = 3'd1;
    assign memory4b[104 ] = 3'd1;
    assign memory4b[105 ] = 3'd1;
    assign memory4b[106 ] = 3'd2;
    assign memory4b[107 ] = 3'd2;
    assign memory4b[108 ] = 3'd2;
    assign memory4b[109 ] = 3'd2;
    assign memory4b[110 ] = 3'd2;
    assign memory4b[111 ] = 3'd2;
    assign memory4b[112 ] = 3'd2;
    assign memory4b[113 ] = 3'd2;
    assign memory4b[114 ] = 3'd2;
    assign memory4b[115 ] = 3'd1;
    assign memory4b[116 ] = 3'd1;
    assign memory4b[117 ] = 3'd1;
    assign memory4b[118 ] = 3'd1;
    assign memory4b[119 ] = 3'd1;
    assign memory4b[120 ] = 3'd2;
    assign memory4b[121 ] = 3'd2;
    assign memory4b[122 ] = 3'd2;
    assign memory4b[123 ] = 3'd2;
    assign memory4b[124 ] = 3'd2;
    assign memory4b[125 ] = 3'd1;
    assign memory4b[126 ] = 3'd1;
    assign memory4b[127 ] = 3'd0;
    assign memory4b[128 ] = 3'd0;
    assign memory4b[129 ] = 3'd1;
    assign memory4b[130 ] = 3'd1;
    assign memory4b[131 ] = 3'd2;
    assign memory4b[132 ] = 3'd2;
    assign memory4b[133 ] = 3'd2;
    assign memory4b[134 ] = 3'd2;
    assign memory4b[135 ] = 3'd2;
    assign memory4b[136 ] = 3'd2;
    assign memory4b[137 ] = 3'd2;
    assign memory4b[138 ] = 3'd2;
    assign memory4b[139 ] = 3'd2;
    assign memory4b[140 ] = 3'd2;
    assign memory4b[141 ] = 3'd2;
    assign memory4b[142 ] = 3'd2;
    assign memory4b[143 ] = 3'd2;
    assign memory4b[144 ] = 3'd2;
    assign memory4b[145 ] = 3'd2;
    assign memory4b[146 ] = 3'd2;
    assign memory4b[147 ] = 3'd2;
    assign memory4b[148 ] = 3'd2;
    assign memory4b[149 ] = 3'd2;
    assign memory4b[150 ] = 3'd2;
    assign memory4b[151 ] = 3'd2;
    assign memory4b[152 ] = 3'd2;
    assign memory4b[153 ] = 3'd2;
    assign memory4b[154 ] = 3'd2;
    assign memory4b[155 ] = 3'd2;
    assign memory4b[156 ] = 3'd2;
    assign memory4b[157 ] = 3'd1;
    assign memory4b[158 ] = 3'd1;
    assign memory4b[159 ] = 3'd0;
    assign memory4b[160 ] = 3'd0;
    assign memory4b[161 ] = 3'd1;
    assign memory4b[162 ] = 3'd1;
    assign memory4b[163 ] = 3'd2;
    assign memory4b[164 ] = 3'd2;
    assign memory4b[165 ] = 3'd2;
    assign memory4b[166 ] = 3'd2;
    assign memory4b[167 ] = 3'd2;
    assign memory4b[168 ] = 3'd2;
    assign memory4b[169 ] = 3'd2;
    assign memory4b[170 ] = 3'd2;
    assign memory4b[171 ] = 3'd2;
    assign memory4b[172 ] = 3'd2;
    assign memory4b[173 ] = 3'd2;
    assign memory4b[174 ] = 3'd2;
    assign memory4b[175 ] = 3'd2;
    assign memory4b[176 ] = 3'd2;
    assign memory4b[177 ] = 3'd2;
    assign memory4b[178 ] = 3'd2;
    assign memory4b[179 ] = 3'd2;
    assign memory4b[180 ] = 3'd2;
    assign memory4b[181 ] = 3'd2;
    assign memory4b[182 ] = 3'd2;
    assign memory4b[183 ] = 3'd2;
    assign memory4b[184 ] = 3'd2;
    assign memory4b[185 ] = 3'd3;
    assign memory4b[186 ] = 3'd2;
    assign memory4b[187 ] = 3'd2;
    assign memory4b[188 ] = 3'd2;
    assign memory4b[189 ] = 3'd1;
    assign memory4b[190 ] = 3'd1;
    assign memory4b[191 ] = 3'd0;
    assign memory4b[192 ] = 3'd0;
    assign memory4b[193 ] = 3'd1;
    assign memory4b[194 ] = 3'd1;
    assign memory4b[195 ] = 3'd1;
    assign memory4b[196 ] = 3'd2;
    assign memory4b[197 ] = 3'd2;
    assign memory4b[198 ] = 3'd2;
    assign memory4b[199 ] = 3'd2;
    assign memory4b[200 ] = 3'd2;
    assign memory4b[201 ] = 3'd2;
    assign memory4b[202 ] = 3'd2;
    assign memory4b[203 ] = 3'd2;
    assign memory4b[204 ] = 3'd2;
    assign memory4b[205 ] = 3'd2;
    assign memory4b[206 ] = 3'd2;
    assign memory4b[207 ] = 3'd2;
    assign memory4b[208 ] = 3'd2;
    assign memory4b[209 ] = 3'd2;
    assign memory4b[210 ] = 3'd2;
    assign memory4b[211 ] = 3'd2;
    assign memory4b[212 ] = 3'd2;
    assign memory4b[213 ] = 3'd2;
    assign memory4b[214 ] = 3'd2;
    assign memory4b[215 ] = 3'd2;
    assign memory4b[216 ] = 3'd2;
    assign memory4b[217 ] = 3'd2;
    assign memory4b[218 ] = 3'd2;
    assign memory4b[219 ] = 3'd2;
    assign memory4b[220 ] = 3'd2;
    assign memory4b[221 ] = 3'd1;
    assign memory4b[222 ] = 3'd1;
    assign memory4b[223 ] = 3'd0;
    assign memory4b[224 ] = 3'd0;
    assign memory4b[225 ] = 3'd1;
    assign memory4b[226 ] = 3'd1;
    assign memory4b[227 ] = 3'd1;
    assign memory4b[228 ] = 3'd2;
    assign memory4b[229 ] = 3'd2;
    assign memory4b[230 ] = 3'd2;
    assign memory4b[231 ] = 3'd2;
    assign memory4b[232 ] = 3'd2;
    assign memory4b[233 ] = 3'd2;
    assign memory4b[234 ] = 3'd3;
    assign memory4b[235 ] = 3'd2;
    assign memory4b[236 ] = 3'd2;
    assign memory4b[237 ] = 3'd2;
    assign memory4b[238 ] = 3'd2;
    assign memory4b[239 ] = 3'd2;
    assign memory4b[240 ] = 3'd2;
    assign memory4b[241 ] = 3'd2;
    assign memory4b[242 ] = 3'd2;
    assign memory4b[243 ] = 3'd2;
    assign memory4b[244 ] = 3'd2;
    assign memory4b[245 ] = 3'd2;
    assign memory4b[246 ] = 3'd2;
    assign memory4b[247 ] = 3'd2;
    assign memory4b[248 ] = 3'd2;
    assign memory4b[249 ] = 3'd2;
    assign memory4b[250 ] = 3'd2;
    assign memory4b[251 ] = 3'd2;
    assign memory4b[252 ] = 3'd2;
    assign memory4b[253 ] = 3'd1;
    assign memory4b[254 ] = 3'd1;
    assign memory4b[255 ] = 3'd0;
    assign memory4b[256 ] = 3'd0;
    assign memory4b[257 ] = 3'd1;
    assign memory4b[258 ] = 3'd1;
    assign memory4b[259 ] = 3'd1;
    assign memory4b[260 ] = 3'd2;
    assign memory4b[261 ] = 3'd2;
    assign memory4b[262 ] = 3'd2;
    assign memory4b[263 ] = 3'd2;
    assign memory4b[264 ] = 3'd2;
    assign memory4b[265 ] = 3'd2;
    assign memory4b[266 ] = 3'd2;
    assign memory4b[267 ] = 3'd2;
    assign memory4b[268 ] = 3'd2;
    assign memory4b[269 ] = 3'd2;
    assign memory4b[270 ] = 3'd2;
    assign memory4b[271 ] = 3'd2;
    assign memory4b[272 ] = 3'd2;
    assign memory4b[273 ] = 3'd2;
    assign memory4b[274 ] = 3'd2;
    assign memory4b[275 ] = 3'd2;
    assign memory4b[276 ] = 3'd3;
    assign memory4b[277 ] = 3'd2;
    assign memory4b[278 ] = 3'd2;
    assign memory4b[279 ] = 3'd2;
    assign memory4b[280 ] = 3'd2;
    assign memory4b[281 ] = 3'd2;
    assign memory4b[282 ] = 3'd2;
    assign memory4b[283 ] = 3'd2;
    assign memory4b[284 ] = 3'd2;
    assign memory4b[285 ] = 3'd1;
    assign memory4b[286 ] = 3'd1;
    assign memory4b[287 ] = 3'd0;
    assign memory4b[288 ] = 3'd0;
    assign memory4b[289 ] = 3'd1;
    assign memory4b[290 ] = 3'd1;
    assign memory4b[291 ] = 3'd2;
    assign memory4b[292 ] = 3'd2;
    assign memory4b[293 ] = 3'd2;
    assign memory4b[294 ] = 3'd2;
    assign memory4b[295 ] = 3'd2;
    assign memory4b[296 ] = 3'd2;
    assign memory4b[297 ] = 3'd2;
    assign memory4b[298 ] = 3'd2;
    assign memory4b[299 ] = 3'd2;
    assign memory4b[300 ] = 3'd2;
    assign memory4b[301 ] = 3'd2;
    assign memory4b[302 ] = 3'd2;
    assign memory4b[303 ] = 3'd2;
    assign memory4b[304 ] = 3'd2;
    assign memory4b[305 ] = 3'd2;
    assign memory4b[306 ] = 3'd2;
    assign memory4b[307 ] = 3'd2;
    assign memory4b[308 ] = 3'd2;
    assign memory4b[309 ] = 3'd2;
    assign memory4b[310 ] = 3'd2;
    assign memory4b[311 ] = 3'd2;
    assign memory4b[312 ] = 3'd2;
    assign memory4b[313 ] = 3'd2;
    assign memory4b[314 ] = 3'd2;
    assign memory4b[315 ] = 3'd2;
    assign memory4b[316 ] = 3'd1;
    assign memory4b[317 ] = 3'd1;
    assign memory4b[318 ] = 3'd1;
    assign memory4b[319 ] = 3'd0;
    assign memory4b[320 ] = 3'd0;
    assign memory4b[321 ] = 3'd1;
    assign memory4b[322 ] = 3'd1;
    assign memory4b[323 ] = 3'd2;
    assign memory4b[324 ] = 3'd2;
    assign memory4b[325 ] = 3'd2;
    assign memory4b[326 ] = 3'd2;
    assign memory4b[327 ] = 3'd2;
    assign memory4b[328 ] = 3'd2;
    assign memory4b[329 ] = 3'd2;
    assign memory4b[330 ] = 3'd2;
    assign memory4b[331 ] = 3'd2;
    assign memory4b[332 ] = 3'd2;
    assign memory4b[333 ] = 3'd2;
    assign memory4b[334 ] = 3'd2;
    assign memory4b[335 ] = 3'd2;
    assign memory4b[336 ] = 3'd2;
    assign memory4b[337 ] = 3'd2;
    assign memory4b[338 ] = 3'd2;
    assign memory4b[339 ] = 3'd2;
    assign memory4b[340 ] = 3'd2;
    assign memory4b[341 ] = 3'd2;
    assign memory4b[342 ] = 3'd2;
    assign memory4b[343 ] = 3'd2;
    assign memory4b[344 ] = 3'd2;
    assign memory4b[345 ] = 3'd2;
    assign memory4b[346 ] = 3'd2;
    assign memory4b[347 ] = 3'd2;
    assign memory4b[348 ] = 3'd1;
    assign memory4b[349 ] = 3'd1;
    assign memory4b[350 ] = 3'd1;
    assign memory4b[351 ] = 3'd0;
    assign memory4b[352 ] = 3'd0;
    assign memory4b[353 ] = 3'd1;
    assign memory4b[354 ] = 3'd1;
    assign memory4b[355 ] = 3'd2;
    assign memory4b[356 ] = 3'd2;
    assign memory4b[357 ] = 3'd2;
    assign memory4b[358 ] = 3'd2;
    assign memory4b[359 ] = 3'd2;
    assign memory4b[360 ] = 3'd2;
    assign memory4b[361 ] = 3'd2;
    assign memory4b[362 ] = 3'd2;
    assign memory4b[363 ] = 3'd2;
    assign memory4b[364 ] = 3'd2;
    assign memory4b[365 ] = 3'd2;
    assign memory4b[366 ] = 3'd2;
    assign memory4b[367 ] = 3'd3;
    assign memory4b[368 ] = 3'd2;
    assign memory4b[369 ] = 3'd2;
    assign memory4b[370 ] = 3'd2;
    assign memory4b[371 ] = 3'd2;
    assign memory4b[372 ] = 3'd2;
    assign memory4b[373 ] = 3'd2;
    assign memory4b[374 ] = 3'd2;
    assign memory4b[375 ] = 3'd2;
    assign memory4b[376 ] = 3'd2;
    assign memory4b[377 ] = 3'd2;
    assign memory4b[378 ] = 3'd2;
    assign memory4b[379 ] = 3'd2;
    assign memory4b[380 ] = 3'd1;
    assign memory4b[381 ] = 3'd1;
    assign memory4b[382 ] = 3'd1;
    assign memory4b[383 ] = 3'd0;
    assign memory4b[384 ] = 3'd0;
    assign memory4b[385 ] = 3'd1;
    assign memory4b[386 ] = 3'd1;
    assign memory4b[387 ] = 3'd2;
    assign memory4b[388 ] = 3'd2;
    assign memory4b[389 ] = 3'd2;
    assign memory4b[390 ] = 3'd2;
    assign memory4b[391 ] = 3'd2;
    assign memory4b[392 ] = 3'd2;
    assign memory4b[393 ] = 3'd2;
    assign memory4b[394 ] = 3'd2;
    assign memory4b[395 ] = 3'd2;
    assign memory4b[396 ] = 3'd2;
    assign memory4b[397 ] = 3'd2;
    assign memory4b[398 ] = 3'd2;
    assign memory4b[399 ] = 3'd2;
    assign memory4b[400 ] = 3'd2;
    assign memory4b[401 ] = 3'd2;
    assign memory4b[402 ] = 3'd2;
    assign memory4b[403 ] = 3'd2;
    assign memory4b[404 ] = 3'd2;
    assign memory4b[405 ] = 3'd2;
    assign memory4b[406 ] = 3'd2;
    assign memory4b[407 ] = 3'd2;
    assign memory4b[408 ] = 3'd2;
    assign memory4b[409 ] = 3'd2;
    assign memory4b[410 ] = 3'd2;
    assign memory4b[411 ] = 3'd2;
    assign memory4b[412 ] = 3'd1;
    assign memory4b[413 ] = 3'd1;
    assign memory4b[414 ] = 3'd1;
    assign memory4b[415 ] = 3'd0;
    assign memory4b[416 ] = 3'd0;
    assign memory4b[417 ] = 3'd1;
    assign memory4b[418 ] = 3'd1;
    assign memory4b[419 ] = 3'd2;
    assign memory4b[420 ] = 3'd2;
    assign memory4b[421 ] = 3'd2;
    assign memory4b[422 ] = 3'd2;
    assign memory4b[423 ] = 3'd2;
    assign memory4b[424 ] = 3'd2;
    assign memory4b[425 ] = 3'd2;
    assign memory4b[426 ] = 3'd2;
    assign memory4b[427 ] = 3'd2;
    assign memory4b[428 ] = 3'd2;
    assign memory4b[429 ] = 3'd2;
    assign memory4b[430 ] = 3'd2;
    assign memory4b[431 ] = 3'd2;
    assign memory4b[432 ] = 3'd2;
    assign memory4b[433 ] = 3'd2;
    assign memory4b[434 ] = 3'd2;
    assign memory4b[435 ] = 3'd2;
    assign memory4b[436 ] = 3'd2;
    assign memory4b[437 ] = 3'd2;
    assign memory4b[438 ] = 3'd2;
    assign memory4b[439 ] = 3'd2;
    assign memory4b[440 ] = 3'd2;
    assign memory4b[441 ] = 3'd2;
    assign memory4b[442 ] = 3'd2;
    assign memory4b[443 ] = 3'd2;
    assign memory4b[444 ] = 3'd1;
    assign memory4b[445 ] = 3'd1;
    assign memory4b[446 ] = 3'd1;
    assign memory4b[447 ] = 3'd0;
    assign memory4b[448 ] = 3'd0;
    assign memory4b[449 ] = 3'd1;
    assign memory4b[450 ] = 3'd1;
    assign memory4b[451 ] = 3'd2;
    assign memory4b[452 ] = 3'd2;
    assign memory4b[453 ] = 3'd2;
    assign memory4b[454 ] = 3'd2;
    assign memory4b[455 ] = 3'd2;
    assign memory4b[456 ] = 3'd3;
    assign memory4b[457 ] = 3'd2;
    assign memory4b[458 ] = 3'd2;
    assign memory4b[459 ] = 3'd2;
    assign memory4b[460 ] = 3'd2;
    assign memory4b[461 ] = 3'd2;
    assign memory4b[462 ] = 3'd3;
    assign memory4b[463 ] = 3'd2;
    assign memory4b[464 ] = 3'd2;
    assign memory4b[465 ] = 3'd2;
    assign memory4b[466 ] = 3'd2;
    assign memory4b[467 ] = 3'd2;
    assign memory4b[468 ] = 3'd2;
    assign memory4b[469 ] = 3'd2;
    assign memory4b[470 ] = 3'd3;
    assign memory4b[471 ] = 3'd2;
    assign memory4b[472 ] = 3'd2;
    assign memory4b[473 ] = 3'd2;
    assign memory4b[474 ] = 3'd2;
    assign memory4b[475 ] = 3'd2;
    assign memory4b[476 ] = 3'd2;
    assign memory4b[477 ] = 3'd1;
    assign memory4b[478 ] = 3'd1;
    assign memory4b[479 ] = 3'd0;
    assign memory4b[480 ] = 3'd0;
    assign memory4b[481 ] = 3'd1;
    assign memory4b[482 ] = 3'd1;
    assign memory4b[483 ] = 3'd2;
    assign memory4b[484 ] = 3'd2;
    assign memory4b[485 ] = 3'd2;
    assign memory4b[486 ] = 3'd2;
    assign memory4b[487 ] = 3'd2;
    assign memory4b[488 ] = 3'd2;
    assign memory4b[489 ] = 3'd2;
    assign memory4b[490 ] = 3'd2;
    assign memory4b[491 ] = 3'd2;
    assign memory4b[492 ] = 3'd2;
    assign memory4b[493 ] = 3'd2;
    assign memory4b[494 ] = 3'd2;
    assign memory4b[495 ] = 3'd2;
    assign memory4b[496 ] = 3'd2;
    assign memory4b[497 ] = 3'd2;
    assign memory4b[498 ] = 3'd2;
    assign memory4b[499 ] = 3'd2;
    assign memory4b[500 ] = 3'd2;
    assign memory4b[501 ] = 3'd2;
    assign memory4b[502 ] = 3'd2;
    assign memory4b[503 ] = 3'd2;
    assign memory4b[504 ] = 3'd2;
    assign memory4b[505 ] = 3'd2;
    assign memory4b[506 ] = 3'd2;
    assign memory4b[507 ] = 3'd2;
    assign memory4b[508 ] = 3'd2;
    assign memory4b[509 ] = 3'd1;
    assign memory4b[510 ] = 3'd1;
    assign memory4b[511 ] = 3'd0;
    assign memory4b[512 ] = 3'd0;
    assign memory4b[513 ] = 3'd1;
    assign memory4b[514 ] = 3'd1;
    assign memory4b[515 ] = 3'd2;
    assign memory4b[516 ] = 3'd2;
    assign memory4b[517 ] = 3'd2;
    assign memory4b[518 ] = 3'd2;
    assign memory4b[519 ] = 3'd2;
    assign memory4b[520 ] = 3'd2;
    assign memory4b[521 ] = 3'd2;
    assign memory4b[522 ] = 3'd2;
    assign memory4b[523 ] = 3'd2;
    assign memory4b[524 ] = 3'd2;
    assign memory4b[525 ] = 3'd2;
    assign memory4b[526 ] = 3'd2;
    assign memory4b[527 ] = 3'd2;
    assign memory4b[528 ] = 3'd2;
    assign memory4b[529 ] = 3'd2;
    assign memory4b[530 ] = 3'd2;
    assign memory4b[531 ] = 3'd2;
    assign memory4b[532 ] = 3'd2;
    assign memory4b[533 ] = 3'd2;
    assign memory4b[534 ] = 3'd2;
    assign memory4b[535 ] = 3'd2;
    assign memory4b[536 ] = 3'd2;
    assign memory4b[537 ] = 3'd2;
    assign memory4b[538 ] = 3'd2;
    assign memory4b[539 ] = 3'd2;
    assign memory4b[540 ] = 3'd2;
    assign memory4b[541 ] = 3'd1;
    assign memory4b[542 ] = 3'd1;
    assign memory4b[543 ] = 3'd0;
    assign memory4b[544 ] = 3'd0;
    assign memory4b[545 ] = 3'd1;
    assign memory4b[546 ] = 3'd1;
    assign memory4b[547 ] = 3'd2;
    assign memory4b[548 ] = 3'd2;
    assign memory4b[549 ] = 3'd2;
    assign memory4b[550 ] = 3'd2;
    assign memory4b[551 ] = 3'd2;
    assign memory4b[552 ] = 3'd2;
    assign memory4b[553 ] = 3'd2;
    assign memory4b[554 ] = 3'd2;
    assign memory4b[555 ] = 3'd2;
    assign memory4b[556 ] = 3'd2;
    assign memory4b[557 ] = 3'd2;
    assign memory4b[558 ] = 3'd2;
    assign memory4b[559 ] = 3'd2;
    assign memory4b[560 ] = 3'd3;
    assign memory4b[561 ] = 3'd2;
    assign memory4b[562 ] = 3'd2;
    assign memory4b[563 ] = 3'd2;
    assign memory4b[564 ] = 3'd2;
    assign memory4b[565 ] = 3'd2;
    assign memory4b[566 ] = 3'd2;
    assign memory4b[567 ] = 3'd2;
    assign memory4b[568 ] = 3'd2;
    assign memory4b[569 ] = 3'd2;
    assign memory4b[570 ] = 3'd2;
    assign memory4b[571 ] = 3'd2;
    assign memory4b[572 ] = 3'd2;
    assign memory4b[573 ] = 3'd1;
    assign memory4b[574 ] = 3'd1;
    assign memory4b[575 ] = 3'd0;
    assign memory4b[576 ] = 3'd0;
    assign memory4b[577 ] = 3'd1;
    assign memory4b[578 ] = 3'd1;
    assign memory4b[579 ] = 3'd2;
    assign memory4b[580 ] = 3'd2;
    assign memory4b[581 ] = 3'd2;
    assign memory4b[582 ] = 3'd2;
    assign memory4b[583 ] = 3'd2;
    assign memory4b[584 ] = 3'd2;
    assign memory4b[585 ] = 3'd2;
    assign memory4b[586 ] = 3'd2;
    assign memory4b[587 ] = 3'd2;
    assign memory4b[588 ] = 3'd2;
    assign memory4b[589 ] = 3'd2;
    assign memory4b[590 ] = 3'd2;
    assign memory4b[591 ] = 3'd2;
    assign memory4b[592 ] = 3'd2;
    assign memory4b[593 ] = 3'd2;
    assign memory4b[594 ] = 3'd2;
    assign memory4b[595 ] = 3'd2;
    assign memory4b[596 ] = 3'd2;
    assign memory4b[597 ] = 3'd2;
    assign memory4b[598 ] = 3'd2;
    assign memory4b[599 ] = 3'd2;
    assign memory4b[600 ] = 3'd2;
    assign memory4b[601 ] = 3'd3;
    assign memory4b[602 ] = 3'd2;
    assign memory4b[603 ] = 3'd2;
    assign memory4b[604 ] = 3'd1;
    assign memory4b[605 ] = 3'd1;
    assign memory4b[606 ] = 3'd1;
    assign memory4b[607 ] = 3'd0;
    assign memory4b[608 ] = 3'd0;
    assign memory4b[609 ] = 3'd1;
    assign memory4b[610 ] = 3'd1;
    assign memory4b[611 ] = 3'd1;
    assign memory4b[612 ] = 3'd2;
    assign memory4b[613 ] = 3'd2;
    assign memory4b[614 ] = 3'd2;
    assign memory4b[615 ] = 3'd2;
    assign memory4b[616 ] = 3'd2;
    assign memory4b[617 ] = 3'd2;
    assign memory4b[618 ] = 3'd2;
    assign memory4b[619 ] = 3'd2;
    assign memory4b[620 ] = 3'd2;
    assign memory4b[621 ] = 3'd2;
    assign memory4b[622 ] = 3'd2;
    assign memory4b[623 ] = 3'd2;
    assign memory4b[624 ] = 3'd2;
    assign memory4b[625 ] = 3'd2;
    assign memory4b[626 ] = 3'd2;
    assign memory4b[627 ] = 3'd2;
    assign memory4b[628 ] = 3'd2;
    assign memory4b[629 ] = 3'd2;
    assign memory4b[630 ] = 3'd2;
    assign memory4b[631 ] = 3'd2;
    assign memory4b[632 ] = 3'd2;
    assign memory4b[633 ] = 3'd3;
    assign memory4b[634 ] = 3'd2;
    assign memory4b[635 ] = 3'd2;
    assign memory4b[636 ] = 3'd1;
    assign memory4b[637 ] = 3'd1;
    assign memory4b[638 ] = 3'd1;
    assign memory4b[639 ] = 3'd0;
    assign memory4b[640 ] = 3'd0;
    assign memory4b[641 ] = 3'd1;
    assign memory4b[642 ] = 3'd1;
    assign memory4b[643 ] = 3'd1;
    assign memory4b[644 ] = 3'd2;
    assign memory4b[645 ] = 3'd2;
    assign memory4b[646 ] = 3'd2;
    assign memory4b[647 ] = 3'd2;
    assign memory4b[648 ] = 3'd2;
    assign memory4b[649 ] = 3'd2;
    assign memory4b[650 ] = 3'd2;
    assign memory4b[651 ] = 3'd2;
    assign memory4b[652 ] = 3'd2;
    assign memory4b[653 ] = 3'd2;
    assign memory4b[654 ] = 3'd2;
    assign memory4b[655 ] = 3'd2;
    assign memory4b[656 ] = 3'd2;
    assign memory4b[657 ] = 3'd2;
    assign memory4b[658 ] = 3'd2;
    assign memory4b[659 ] = 3'd2;
    assign memory4b[660 ] = 3'd2;
    assign memory4b[661 ] = 3'd2;
    assign memory4b[662 ] = 3'd2;
    assign memory4b[663 ] = 3'd2;
    assign memory4b[664 ] = 3'd2;
    assign memory4b[665 ] = 3'd2;
    assign memory4b[666 ] = 3'd2;
    assign memory4b[667 ] = 3'd2;
    assign memory4b[668 ] = 3'd1;
    assign memory4b[669 ] = 3'd1;
    assign memory4b[670 ] = 3'd1;
    assign memory4b[671 ] = 3'd0;
    assign memory4b[672 ] = 3'd0;
    assign memory4b[673 ] = 3'd1;
    assign memory4b[674 ] = 3'd1;
    assign memory4b[675 ] = 3'd1;
    assign memory4b[676 ] = 3'd2;
    assign memory4b[677 ] = 3'd2;
    assign memory4b[678 ] = 3'd2;
    assign memory4b[679 ] = 3'd2;
    assign memory4b[680 ] = 3'd2;
    assign memory4b[681 ] = 3'd2;
    assign memory4b[682 ] = 3'd2;
    assign memory4b[683 ] = 3'd2;
    assign memory4b[684 ] = 3'd2;
    assign memory4b[685 ] = 3'd2;
    assign memory4b[686 ] = 3'd2;
    assign memory4b[687 ] = 3'd2;
    assign memory4b[688 ] = 3'd2;
    assign memory4b[689 ] = 3'd2;
    assign memory4b[690 ] = 3'd2;
    assign memory4b[691 ] = 3'd2;
    assign memory4b[692 ] = 3'd2;
    assign memory4b[693 ] = 3'd2;
    assign memory4b[694 ] = 3'd2;
    assign memory4b[695 ] = 3'd2;
    assign memory4b[696 ] = 3'd2;
    assign memory4b[697 ] = 3'd2;
    assign memory4b[698 ] = 3'd2;
    assign memory4b[699 ] = 3'd2;
    assign memory4b[700 ] = 3'd1;
    assign memory4b[701 ] = 3'd1;
    assign memory4b[702 ] = 3'd1;
    assign memory4b[703 ] = 3'd0;
    assign memory4b[704 ] = 3'd0;
    assign memory4b[705 ] = 3'd1;
    assign memory4b[706 ] = 3'd1;
    assign memory4b[707 ] = 3'd1;
    assign memory4b[708 ] = 3'd2;
    assign memory4b[709 ] = 3'd2;
    assign memory4b[710 ] = 3'd2;
    assign memory4b[711 ] = 3'd2;
    assign memory4b[712 ] = 3'd2;
    assign memory4b[713 ] = 3'd2;
    assign memory4b[714 ] = 3'd2;
    assign memory4b[715 ] = 3'd2;
    assign memory4b[716 ] = 3'd2;
    assign memory4b[717 ] = 3'd3;
    assign memory4b[718 ] = 3'd2;
    assign memory4b[719 ] = 3'd2;
    assign memory4b[720 ] = 3'd2;
    assign memory4b[721 ] = 3'd2;
    assign memory4b[722 ] = 3'd2;
    assign memory4b[723 ] = 3'd2;
    assign memory4b[724 ] = 3'd2;
    assign memory4b[725 ] = 3'd2;
    assign memory4b[726 ] = 3'd2;
    assign memory4b[727 ] = 3'd2;
    assign memory4b[728 ] = 3'd2;
    assign memory4b[729 ] = 3'd2;
    assign memory4b[730 ] = 3'd2;
    assign memory4b[731 ] = 3'd2;
    assign memory4b[732 ] = 3'd2;
    assign memory4b[733 ] = 3'd1;
    assign memory4b[734 ] = 3'd1;
    assign memory4b[735 ] = 3'd0;
    assign memory4b[736 ] = 3'd0;
    assign memory4b[737 ] = 3'd1;
    assign memory4b[738 ] = 3'd1;
    assign memory4b[739 ] = 3'd1;
    assign memory4b[740 ] = 3'd2;
    assign memory4b[741 ] = 3'd2;
    assign memory4b[742 ] = 3'd2;
    assign memory4b[743 ] = 3'd2;
    assign memory4b[744 ] = 3'd3;
    assign memory4b[745 ] = 3'd2;
    assign memory4b[746 ] = 3'd2;
    assign memory4b[747 ] = 3'd2;
    assign memory4b[748 ] = 3'd2;
    assign memory4b[749 ] = 3'd2;
    assign memory4b[750 ] = 3'd2;
    assign memory4b[751 ] = 3'd2;
    assign memory4b[752 ] = 3'd2;
    assign memory4b[753 ] = 3'd2;
    assign memory4b[754 ] = 3'd2;
    assign memory4b[755 ] = 3'd2;
    assign memory4b[756 ] = 3'd2;
    assign memory4b[757 ] = 3'd2;
    assign memory4b[758 ] = 3'd3;
    assign memory4b[759 ] = 3'd2;
    assign memory4b[760 ] = 3'd2;
    assign memory4b[761 ] = 3'd2;
    assign memory4b[762 ] = 3'd2;
    assign memory4b[763 ] = 3'd2;
    assign memory4b[764 ] = 3'd2;
    assign memory4b[765 ] = 3'd1;
    assign memory4b[766 ] = 3'd1;
    assign memory4b[767 ] = 3'd0;
    assign memory4b[768 ] = 3'd0;
    assign memory4b[769 ] = 3'd1;
    assign memory4b[770 ] = 3'd1;
    assign memory4b[771 ] = 3'd2;
    assign memory4b[772 ] = 3'd2;
    assign memory4b[773 ] = 3'd2;
    assign memory4b[774 ] = 3'd2;
    assign memory4b[775 ] = 3'd2;
    assign memory4b[776 ] = 3'd2;
    assign memory4b[777 ] = 3'd2;
    assign memory4b[778 ] = 3'd2;
    assign memory4b[779 ] = 3'd2;
    assign memory4b[780 ] = 3'd2;
    assign memory4b[781 ] = 3'd2;
    assign memory4b[782 ] = 3'd2;
    assign memory4b[783 ] = 3'd2;
    assign memory4b[784 ] = 3'd2;
    assign memory4b[785 ] = 3'd2;
    assign memory4b[786 ] = 3'd2;
    assign memory4b[787 ] = 3'd2;
    assign memory4b[788 ] = 3'd2;
    assign memory4b[789 ] = 3'd2;
    assign memory4b[790 ] = 3'd2;
    assign memory4b[791 ] = 3'd2;
    assign memory4b[792 ] = 3'd2;
    assign memory4b[793 ] = 3'd2;
    assign memory4b[794 ] = 3'd2;
    assign memory4b[795 ] = 3'd2;
    assign memory4b[796 ] = 3'd2;
    assign memory4b[797 ] = 3'd1;
    assign memory4b[798 ] = 3'd1;
    assign memory4b[799 ] = 3'd0;
    assign memory4b[800 ] = 3'd0;
    assign memory4b[801 ] = 3'd1;
    assign memory4b[802 ] = 3'd1;
    assign memory4b[803 ] = 3'd2;
    assign memory4b[804 ] = 3'd2;
    assign memory4b[805 ] = 3'd2;
    assign memory4b[806 ] = 3'd2;
    assign memory4b[807 ] = 3'd2;
    assign memory4b[808 ] = 3'd2;
    assign memory4b[809 ] = 3'd2;
    assign memory4b[810 ] = 3'd2;
    assign memory4b[811 ] = 3'd2;
    assign memory4b[812 ] = 3'd2;
    assign memory4b[813 ] = 3'd2;
    assign memory4b[814 ] = 3'd2;
    assign memory4b[815 ] = 3'd2;
    assign memory4b[816 ] = 3'd2;
    assign memory4b[817 ] = 3'd2;
    assign memory4b[818 ] = 3'd2;
    assign memory4b[819 ] = 3'd2;
    assign memory4b[820 ] = 3'd2;
    assign memory4b[821 ] = 3'd2;
    assign memory4b[822 ] = 3'd2;
    assign memory4b[823 ] = 3'd2;
    assign memory4b[824 ] = 3'd2;
    assign memory4b[825 ] = 3'd2;
    assign memory4b[826 ] = 3'd3;
    assign memory4b[827 ] = 3'd2;
    assign memory4b[828 ] = 3'd2;
    assign memory4b[829 ] = 3'd1;
    assign memory4b[830 ] = 3'd1;
    assign memory4b[831 ] = 3'd0;
    assign memory4b[832 ] = 3'd0;
    assign memory4b[833 ] = 3'd1;
    assign memory4b[834 ] = 3'd1;
    assign memory4b[835 ] = 3'd2;
    assign memory4b[836 ] = 3'd2;
    assign memory4b[837 ] = 3'd2;
    assign memory4b[838 ] = 3'd2;
    assign memory4b[839 ] = 3'd2;
    assign memory4b[840 ] = 3'd2;
    assign memory4b[841 ] = 3'd2;
    assign memory4b[842 ] = 3'd2;
    assign memory4b[843 ] = 3'd2;
    assign memory4b[844 ] = 3'd2;
    assign memory4b[845 ] = 3'd2;
    assign memory4b[846 ] = 3'd2;
    assign memory4b[847 ] = 3'd2;
    assign memory4b[848 ] = 3'd2;
    assign memory4b[849 ] = 3'd2;
    assign memory4b[850 ] = 3'd2;
    assign memory4b[851 ] = 3'd2;
    assign memory4b[852 ] = 3'd2;
    assign memory4b[853 ] = 3'd2;
    assign memory4b[854 ] = 3'd2;
    assign memory4b[855 ] = 3'd2;
    assign memory4b[856 ] = 3'd2;
    assign memory4b[857 ] = 3'd2;
    assign memory4b[858 ] = 3'd2;
    assign memory4b[859 ] = 3'd2;
    assign memory4b[860 ] = 3'd1;
    assign memory4b[861 ] = 3'd1;
    assign memory4b[862 ] = 3'd1;
    assign memory4b[863 ] = 3'd0;
    assign memory4b[864 ] = 3'd0;
    assign memory4b[865 ] = 3'd1;
    assign memory4b[866 ] = 3'd1;
    assign memory4b[867 ] = 3'd2;
    assign memory4b[868 ] = 3'd2;
    assign memory4b[869 ] = 3'd2;
    assign memory4b[870 ] = 3'd2;
    assign memory4b[871 ] = 3'd2;
    assign memory4b[872 ] = 3'd2;
    assign memory4b[873 ] = 3'd2;
    assign memory4b[874 ] = 3'd2;
    assign memory4b[875 ] = 3'd2;
    assign memory4b[876 ] = 3'd2;
    assign memory4b[877 ] = 3'd2;
    assign memory4b[878 ] = 3'd2;
    assign memory4b[879 ] = 3'd2;
    assign memory4b[880 ] = 3'd2;
    assign memory4b[881 ] = 3'd2;
    assign memory4b[882 ] = 3'd2;
    assign memory4b[883 ] = 3'd2;
    assign memory4b[884 ] = 3'd2;
    assign memory4b[885 ] = 3'd2;
    assign memory4b[886 ] = 3'd2;
    assign memory4b[887 ] = 3'd2;
    assign memory4b[888 ] = 3'd2;
    assign memory4b[889 ] = 3'd2;
    assign memory4b[890 ] = 3'd2;
    assign memory4b[891 ] = 3'd2;
    assign memory4b[892 ] = 3'd1;
    assign memory4b[893 ] = 3'd1;
    assign memory4b[894 ] = 3'd1;
    assign memory4b[895 ] = 3'd0;
    assign memory4b[896 ] = 3'd0;
    assign memory4b[897 ] = 3'd1;
    assign memory4b[898 ] = 3'd1;
    assign memory4b[899 ] = 3'd2;
    assign memory4b[900 ] = 3'd2;
    assign memory4b[901 ] = 3'd2;
    assign memory4b[902 ] = 3'd2;
    assign memory4b[903 ] = 3'd1;
    assign memory4b[904 ] = 3'd1;
    assign memory4b[905 ] = 3'd1;
    assign memory4b[906 ] = 3'd1;
    assign memory4b[907 ] = 3'd2;
    assign memory4b[908 ] = 3'd2;
    assign memory4b[909 ] = 3'd2;
    assign memory4b[910 ] = 3'd1;
    assign memory4b[911 ] = 3'd1;
    assign memory4b[912 ] = 3'd1;
    assign memory4b[913 ] = 3'd2;
    assign memory4b[914 ] = 3'd2;
    assign memory4b[915 ] = 3'd2;
    assign memory4b[916 ] = 3'd2;
    assign memory4b[917 ] = 3'd1;
    assign memory4b[918 ] = 3'd1;
    assign memory4b[919 ] = 3'd1;
    assign memory4b[920 ] = 3'd2;
    assign memory4b[921 ] = 3'd2;
    assign memory4b[922 ] = 3'd2;
    assign memory4b[923 ] = 3'd2;
    assign memory4b[924 ] = 3'd2;
    assign memory4b[925 ] = 3'd1;
    assign memory4b[926 ] = 3'd1;
    assign memory4b[927 ] = 3'd0;
    assign memory4b[928 ] = 3'd0;
    assign memory4b[929 ] = 3'd1;
    assign memory4b[930 ] = 3'd1;
    assign memory4b[931 ] = 3'd1;
    assign memory4b[932 ] = 3'd1;
    assign memory4b[933 ] = 3'd1;
    assign memory4b[934 ] = 3'd1;
    assign memory4b[935 ] = 3'd1;
    assign memory4b[936 ] = 3'd1;
    assign memory4b[937 ] = 3'd1;
    assign memory4b[938 ] = 3'd1;
    assign memory4b[939 ] = 3'd1;
    assign memory4b[940 ] = 3'd1;
    assign memory4b[941 ] = 3'd1;
    assign memory4b[942 ] = 3'd1;
    assign memory4b[943 ] = 3'd1;
    assign memory4b[944 ] = 3'd1;
    assign memory4b[945 ] = 3'd1;
    assign memory4b[946 ] = 3'd1;
    assign memory4b[947 ] = 3'd1;
    assign memory4b[948 ] = 3'd1;
    assign memory4b[949 ] = 3'd1;
    assign memory4b[950 ] = 3'd1;
    assign memory4b[951 ] = 3'd1;
    assign memory4b[952 ] = 3'd1;
    assign memory4b[953 ] = 3'd1;
    assign memory4b[954 ] = 3'd1;
    assign memory4b[955 ] = 3'd1;
    assign memory4b[956 ] = 3'd1;
    assign memory4b[957 ] = 3'd1;
    assign memory4b[958 ] = 3'd1;
    assign memory4b[959 ] = 3'd0;
    assign memory4b[960 ] = 3'd0;
    assign memory4b[961 ] = 3'd1;
    assign memory4b[962 ] = 3'd1;
    assign memory4b[963 ] = 3'd1;
    assign memory4b[964 ] = 3'd1;
    assign memory4b[965 ] = 3'd1;
    assign memory4b[966 ] = 3'd1;
    assign memory4b[967 ] = 3'd1;
    assign memory4b[968 ] = 3'd1;
    assign memory4b[969 ] = 3'd1;
    assign memory4b[970 ] = 3'd1;
    assign memory4b[971 ] = 3'd1;
    assign memory4b[972 ] = 3'd1;
    assign memory4b[973 ] = 3'd1;
    assign memory4b[974 ] = 3'd1;
    assign memory4b[975 ] = 3'd1;
    assign memory4b[976 ] = 3'd1;
    assign memory4b[977 ] = 3'd1;
    assign memory4b[978 ] = 3'd1;
    assign memory4b[979 ] = 3'd1;
    assign memory4b[980 ] = 3'd1;
    assign memory4b[981 ] = 3'd1;
    assign memory4b[982 ] = 3'd1;
    assign memory4b[983 ] = 3'd1;
    assign memory4b[984 ] = 3'd1;
    assign memory4b[985 ] = 3'd1;
    assign memory4b[986 ] = 3'd1;
    assign memory4b[987 ] = 3'd1;
    assign memory4b[988 ] = 3'd1;
    assign memory4b[989 ] = 3'd1;
    assign memory4b[990 ] = 3'd1;
    assign memory4b[991 ] = 3'd0;
    assign memory4b[992 ] = 3'd0;
    assign memory4b[993 ] = 3'd0;
    assign memory4b[994 ] = 3'd0;
    assign memory4b[995 ] = 3'd0;
    assign memory4b[996 ] = 3'd0;
    assign memory4b[997 ] = 3'd0;
    assign memory4b[998 ] = 3'd0;
    assign memory4b[999 ] = 3'd0;
    assign memory4b[1000] = 3'd0;
    assign memory4b[1001] = 3'd0;
    assign memory4b[1002] = 3'd0;
    assign memory4b[1003] = 3'd0;
    assign memory4b[1004] = 3'd0;
    assign memory4b[1005] = 3'd0;
    assign memory4b[1006] = 3'd0;
    assign memory4b[1007] = 3'd0;
    assign memory4b[1008] = 3'd0;
    assign memory4b[1009] = 3'd0;
    assign memory4b[1010] = 3'd0;
    assign memory4b[1011] = 3'd0;
    assign memory4b[1012] = 3'd0;
    assign memory4b[1013] = 3'd0;
    assign memory4b[1014] = 3'd0;
    assign memory4b[1015] = 3'd0;
    assign memory4b[1016] = 3'd0;
    assign memory4b[1017] = 3'd0;
    assign memory4b[1018] = 3'd0;
    assign memory4b[1019] = 3'd0;
    assign memory4b[1020] = 3'd0;
    assign memory4b[1021] = 3'd0;
    assign memory4b[1022] = 3'd0;
    assign memory4b[1023] = 3'd0;

endmodule
