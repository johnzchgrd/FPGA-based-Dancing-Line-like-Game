//	How to use:	
//	1. Edit the songs on the Enter Song sheet.	
// 	2. Select this whole worksheet, copy it, and paste it into a new file.	
//	3. Save the file as song_rom.v.	

module pulse4_rom (
    input clk,						
	output reg [25:0] dout,						
	input [11:0] addr		
    );
        
    wire [25:0] memory [4095:0];        				
	always @(posedge clk)						
		dout = memory[addr];					

    parameter s1 = 402;
    parameter s2 = s1 + 120;
    parameter s3 = s2 + 125;

    assign memory[0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[43 ] = {7'd0  , 8'd234, 7'd0  , 2'd0, 2'd0};
    assign memory[44 ] = {7'd69 , 8'd24 , 7'd92 , 2'd3, 2'd0};   //note: 7F
    assign memory[45 ] = {7'd66 , 8'd24 , 7'd92 , 2'd3, 2'd0};   //note: 7D
    assign memory[46 ] = {7'd64 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 7C
    assign memory[47 ] = {7'd61 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[48 ] = {7'd59 , 8'd32 , 7'd94 , 2'd3, 2'd0};   //note: 6G
    assign memory[49 ] = {7'd57 , 8'd32 , 7'd94 , 2'd3, 2'd0};   //note: 6F
    assign memory[50 ] = {7'd56 , 8'd32 , 7'd94 , 2'd3, 2'd0};   //note: 6E
    assign memory[51 ] = {7'd54 , 8'd4  , 7'd96 , 2'd3, 2'd0};   //note: 6D
    assign memory[52 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[53 ] = {7'd54 , 8'd4  , 7'd96 , 2'd3, 2'd0};   //note: 6D
    assign memory[54 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[55 ] = {7'd54 , 8'd4  , 7'd96 , 2'd3, 2'd0};   //note: 6D
    assign memory[56 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[57 ] = {7'd54 , 8'd4  , 7'd73 , 2'd3, 2'd0};   //note: 6D
    assign memory[58 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[59 ] = {7'd54 , 8'd4  , 7'd62 , 2'd3, 2'd0};   //note: 6D
    assign memory[60 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[61 ] = {7'd54 , 8'd4  , 7'd98 , 2'd3, 2'd0};   //note: 6D
    assign memory[62 ] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[63 ] = {7'd54 , 8'd4  , 7'd98 , 2'd3, 2'd0};   //note: 6D
    assign memory[64 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[65 ] = {7'd54 , 8'd4  , 7'd98 , 2'd3, 2'd0};   //note: 6D
    assign memory[66 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[67 ] = {7'd54 , 8'd4  , 7'd98 , 2'd3, 2'd0};   //note: 6D
    assign memory[68 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[69 ] = {7'd54 , 8'd4  , 7'd98 , 2'd3, 2'd0};   //note: 6D
    assign memory[70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[71 ] = {7'd0  , 8'd246, 7'd0  , 2'd0, 2'd0};
    assign memory[72 ] = {7'd57 , 8'd23 , 7'd100, 2'd3, 2'd0};   //note: 6F
    assign memory[73 ] = {7'd52 , 8'd24 , 7'd101, 2'd3, 2'd0};   //note: 6C
    assign memory[74 ] = {7'd54 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 6D
    assign memory[75 ] = {7'd57 , 8'd24 , 7'd100, 2'd3, 2'd0};   //note: 6F
    assign memory[76 ] = {7'd59 , 8'd23 , 7'd103, 2'd3, 2'd0};   //note: 6G
    assign memory[77 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[78 ] = {7'd57 , 8'd24 , 7'd100, 2'd3, 2'd0};   //note: 6F
    assign memory[79 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[80 ] = {7'd59 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 6G
    assign memory[81 ] = {7'd0  , 8'd10 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[82 ] = {7'd61 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[83 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[84 ] = {7'd61 , 8'd4  , 7'd100, 2'd3, 2'd0};   //note: 6A
    assign memory[85 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[86 ] = {7'd61 , 8'd4  , 7'd100, 2'd3, 2'd0};   //note: 6A
    assign memory[87 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[88 ] = {7'd61 , 8'd4  , 7'd100, 2'd3, 2'd0};   //note: 6A
    assign memory[89 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[90 ] = {7'd61 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[91 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[92 ] = {7'd61 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[93 ] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[94 ] = {7'd61 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[95 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[96 ] = {7'd61 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[97 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[98 ] = {7'd61 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[99 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[100] = {7'd61 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[101] = {7'd0  , 8'd117, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[102] = {7'd64 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 7C
    assign memory[103] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[104] = {7'd61 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[105] = {7'd64 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 7C
    assign memory[106] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[107] = {7'd61 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[108] = {7'd64 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 7C
    assign memory[109] = {7'd0  , 8'd216, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[110] = {7'd69 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 7F
    assign memory[111] = {7'd66 , 8'd24 , 7'd101, 2'd3, 2'd0};   //note: 7D
    assign memory[112] = {7'd64 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 7C
    assign memory[113] = {7'd61 , 8'd24 , 7'd103, 2'd3, 2'd0};   //note: 6A
    assign memory[114] = {7'd59 , 8'd32 , 7'd103, 2'd3, 2'd0};   //note: 6G
    assign memory[115] = {7'd57 , 8'd32 , 7'd103, 2'd3, 2'd0};   //note: 6F
    assign memory[116] = {7'd56 , 8'd32 , 7'd103, 2'd3, 2'd0};   //note: 6E
    assign memory[117] = {7'd54 , 8'd4  , 7'd101, 2'd3, 2'd0};   //note: 6D
    assign memory[118] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[119] = {7'd54 , 8'd4  , 7'd101, 2'd3, 2'd0};   //note: 6D
    assign memory[120] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[121] = {7'd54 , 8'd4  , 7'd84 , 2'd3, 2'd0};   //note: 6D
    assign memory[122] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[123] = {7'd54 , 8'd4  , 7'd73 , 2'd3, 2'd0};   //note: 6D
    assign memory[124] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[125] = {7'd54 , 8'd4  , 7'd62 , 2'd3, 2'd0};   //note: 6D
    assign memory[126] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[127] = {7'd54 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6D
    assign memory[128] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[129] = {7'd54 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6D
    assign memory[130] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[131] = {7'd54 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6D
    assign memory[132] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[133] = {7'd54 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6D
    assign memory[134] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[135] = {7'd54 , 8'd4  , 7'd103, 2'd3, 2'd0};   //note: 6D
    assign memory[136] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[137] = {7'd0  , 8'd246, 7'd0  , 2'd0, 2'd0};
    assign memory[138] = {7'd57 , 8'd23 , 7'd108, 2'd3, 2'd0};   //note: 6F
    assign memory[139] = {7'd52 , 8'd24 , 7'd108, 2'd3, 2'd0};   //note: 6C
    assign memory[140] = {7'd54 , 8'd24 , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[141] = {7'd57 , 8'd24 , 7'd108, 2'd3, 2'd0};   //note: 6F
    assign memory[142] = {7'd59 , 8'd23 , 7'd108, 2'd3, 2'd0};   //note: 6G
    assign memory[143] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[144] = {7'd57 , 8'd24 , 7'd108, 2'd3, 2'd0};   //note: 6F
    assign memory[145] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[146] = {7'd59 , 8'd24 , 7'd108, 2'd3, 2'd0};   //note: 6G
    assign memory[147] = {7'd0  , 8'd10 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[148] = {7'd61 , 8'd4  , 7'd108, 2'd3, 2'd0};   //note: 6A
    assign memory[149] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[150] = {7'd61 , 8'd4  , 7'd108, 2'd3, 2'd0};   //note: 6A
    assign memory[151] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[152] = {7'd61 , 8'd4  , 7'd108, 2'd3, 2'd0};   //note: 6A
    assign memory[153] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[154] = {7'd61 , 8'd4  , 7'd101, 2'd3, 2'd0};   //note: 6A
    assign memory[155] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[156] = {7'd61 , 8'd4  , 7'd101, 2'd3, 2'd0};   //note: 6A
    assign memory[157] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[158] = {7'd61 , 8'd4  , 7'd101, 2'd3, 2'd0};   //note: 6A
    assign memory[159] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[160] = {7'd61 , 8'd4  , 7'd41 , 2'd3, 2'd0};   //note: 6A
    assign memory[161] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[162] = {7'd61 , 8'd4  , 7'd31 , 2'd3, 2'd0};   //note: 6A
    assign memory[163] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[164] = {7'd61 , 8'd4  , 7'd108, 2'd3, 2'd0};   //note: 6A
    assign memory[165] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[166] = {7'd61 , 8'd4  , 7'd108, 2'd3, 2'd0};   //note: 6A
    assign memory[167] = {7'd0  , 8'd117, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[168] = {7'd64 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 7C
    assign memory[169] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[170] = {7'd61 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 6A
    assign memory[171] = {7'd64 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 7C
    assign memory[172] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[173] = {7'd61 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 6A
    assign memory[174] = {7'd64 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 7C
    assign memory[175] = {7'd0  , 8'd216, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[176] = {7'd69 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 7F
    assign memory[177] = {7'd66 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 7D
    assign memory[178] = {7'd64 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 7C
    assign memory[179] = {7'd61 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 6A
    assign memory[180] = {7'd59 , 8'd32 , 7'd107, 2'd3, 2'd0};   //note: 6G
    assign memory[181] = {7'd57 , 8'd32 , 7'd98 , 2'd3, 2'd0};   //note: 6F
    assign memory[182] = {7'd56 , 8'd32 , 7'd107, 2'd3, 2'd0};   //note: 6E
    assign memory[183] = {7'd54 , 8'd4  , 7'd99 , 2'd3, 2'd0};   //note: 6D
    assign memory[184] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[185] = {7'd54 , 8'd4  , 7'd94 , 2'd3, 2'd0};   //note: 6D
    assign memory[186] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[187] = {7'd54 , 8'd4  , 7'd98 , 2'd3, 2'd0};   //note: 6D
    assign memory[188] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[189] = {7'd54 , 8'd4  , 7'd98 , 2'd3, 2'd0};   //note: 6D
    assign memory[190] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[191] = {7'd54 , 8'd4  , 7'd98 , 2'd3, 2'd0};   //note: 6D
    assign memory[192] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[193] = {7'd54 , 8'd4  , 7'd110, 2'd3, 2'd0};   //note: 6D
    assign memory[194] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[195] = {7'd54 , 8'd4  , 7'd110, 2'd3, 2'd0};   //note: 6D
    assign memory[196] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[197] = {7'd54 , 8'd4  , 7'd110, 2'd3, 2'd0};   //note: 6D
    assign memory[198] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[199] = {7'd54 , 8'd4  , 7'd110, 2'd3, 2'd0};   //note: 6D
    assign memory[200] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[201] = {7'd54 , 8'd4  , 7'd110, 2'd3, 2'd0};   //note: 6D
    assign memory[202] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[203] = {7'd0  , 8'd246, 7'd0  , 2'd0, 2'd0};
    assign memory[204] = {7'd57 , 8'd23 , 7'd112, 2'd3, 2'd0};   //note: 6F
    assign memory[205] = {7'd52 , 8'd24 , 7'd116, 2'd3, 2'd0};   //note: 6C
    assign memory[206] = {7'd54 , 8'd24 , 7'd92 , 2'd3, 2'd0};   //note: 6D
    assign memory[207] = {7'd57 , 8'd24 , 7'd114, 2'd3, 2'd0};   //note: 6F
    assign memory[208] = {7'd59 , 8'd23 , 7'd114, 2'd3, 2'd0};   //note: 6G
    assign memory[209] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[210] = {7'd57 , 8'd24 , 7'd114, 2'd3, 2'd0};   //note: 6F
    assign memory[211] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[212] = {7'd59 , 8'd24 , 7'd114, 2'd3, 2'd0};   //note: 6G
    assign memory[213] = {7'd0  , 8'd10 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[214] = {7'd61 , 8'd4  , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[215] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[216] = {7'd61 , 8'd4  , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[217] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[218] = {7'd61 , 8'd4  , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[219] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[220] = {7'd61 , 8'd4  , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[221] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[222] = {7'd61 , 8'd4  , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[223] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[224] = {7'd61 , 8'd4  , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[225] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[226] = {7'd61 , 8'd4  , 7'd92 , 2'd3, 2'd0};   //note: 6A
    assign memory[227] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[228] = {7'd61 , 8'd4  , 7'd92 , 2'd3, 2'd0};   //note: 6A
    assign memory[229] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[230] = {7'd61 , 8'd4  , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[231] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[232] = {7'd61 , 8'd4  , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[233] = {7'd0  , 8'd117, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[234] = {7'd64 , 8'd24 , 7'd114, 2'd3, 2'd0};   //note: 7C
    assign memory[235] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[236] = {7'd61 , 8'd24 , 7'd114, 2'd3, 2'd0};   //note: 6A
    assign memory[237] = {7'd64 , 8'd24 , 7'd112, 2'd3, 2'd0};   //note: 7C
    assign memory[238] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[239] = {7'd61 , 8'd24 , 7'd110, 2'd3, 2'd0};   //note: 6A
    assign memory[240] = {7'd64 , 8'd24 , 7'd110, 2'd3, 2'd0};   //note: 7C
    assign memory[241] = {7'd0  , 8'd216, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[242] = {7'd69 , 8'd24 , 7'd107, 2'd3, 2'd0};   //note: 7F
    assign memory[243] = {7'd66 , 8'd24 , 7'd101, 2'd3, 2'd0};   //note: 7D
    assign memory[244] = {7'd64 , 8'd24 , 7'd101, 2'd3, 2'd0};   //note: 7C
    assign memory[245] = {7'd61 , 8'd24 , 7'd101, 2'd3, 2'd0};   //note: 6A
    assign memory[246] = {7'd59 , 8'd32 , 7'd92 , 2'd3, 2'd0};   //note: 6G
    assign memory[247] = {7'd57 , 8'd32 , 7'd101, 2'd3, 2'd0};   //note: 6F
    assign memory[248] = {7'd56 , 8'd32 , 7'd92 , 2'd3, 2'd0};   //note: 6E
    assign memory[249] = {7'd54 , 8'd4  , 7'd101, 2'd3, 2'd0};   //note: 6D
    assign memory[250] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[251] = {7'd54 , 8'd4  , 7'd101, 2'd3, 2'd0};   //note: 6D
    assign memory[252] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[253] = {7'd54 , 8'd4  , 7'd92 , 2'd3, 2'd0};   //note: 6D
    assign memory[254] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[255] = {7'd54 , 8'd4  , 7'd92 , 2'd3, 2'd0};   //note: 6D
    assign memory[256] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[257] = {7'd54 , 8'd4  , 7'd92 , 2'd3, 2'd0};   //note: 6D
    assign memory[258] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[259] = {7'd54 , 8'd4  , 7'd92 , 2'd3, 2'd0};   //note: 6D
    assign memory[260] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[261] = {7'd54 , 8'd4  , 7'd92 , 2'd3, 2'd0};   //note: 6D
    assign memory[262] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[263] = {7'd54 , 8'd4  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[264] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[265] = {7'd54 , 8'd4  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[266] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[267] = {7'd54 , 8'd4  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[268] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[269] = {7'd0  , 8'd246, 7'd0  , 2'd0, 2'd0};
    assign memory[270] = {7'd57 , 8'd23 , 7'd98 , 2'd3, 2'd0};   //note: 6F
    assign memory[271] = {7'd52 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 6C
    assign memory[272] = {7'd54 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 6D
    assign memory[273] = {7'd57 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 6F
    assign memory[274] = {7'd59 , 8'd23 , 7'd94 , 2'd3, 2'd0};   //note: 6G
    assign memory[275] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[276] = {7'd57 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 6F
    assign memory[277] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[278] = {7'd59 , 8'd24 , 7'd89 , 2'd3, 2'd0};   //note: 6G
    assign memory[279] = {7'd0  , 8'd10 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[280] = {7'd61 , 8'd4  , 7'd96 , 2'd3, 2'd0};   //note: 6A
    assign memory[281] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[282] = {7'd61 , 8'd4  , 7'd96 , 2'd3, 2'd0};   //note: 6A
    assign memory[283] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[284] = {7'd61 , 8'd4  , 7'd96 , 2'd3, 2'd0};   //note: 6A
    assign memory[285] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[286] = {7'd61 , 8'd4  , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[287] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[288] = {7'd61 , 8'd4  , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[289] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[290] = {7'd61 , 8'd4  , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[291] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[292] = {7'd61 , 8'd4  , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[293] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[294] = {7'd61 , 8'd4  , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[295] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[296] = {7'd61 , 8'd4  , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[297] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[298] = {7'd61 , 8'd4  , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[299] = {7'd0  , 8'd117, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[300] = {7'd64 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 7C
    assign memory[301] = {7'd61 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 6A
    assign memory[302] = {7'd64 , 8'd48 , 7'd92 , 2'd3, 2'd0};   //note: 7C
    assign memory[303] = {7'd61 , 8'd24 , 7'd92 , 2'd3, 2'd0};   //note: 6A
    assign memory[304] = {7'd64 , 8'd24 , 7'd92 , 2'd3, 2'd0};   //note: 7C
    assign memory[305] = {7'd66 , 8'd24 , 7'd92 , 2'd3, 2'd0};   //note: 7D
    assign memory[306] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[307] = {7'd69 , 8'd8  , 7'd94 , 2'd3, 2'd0};   //note: 7F
    assign memory[308] = {7'd66 , 8'd8  , 7'd92 , 2'd3, 2'd0};   //note: 7D
    assign memory[309] = {7'd69 , 8'd8  , 7'd92 , 2'd3, 2'd0};   //note: 7F
    assign memory[310] = {7'd66 , 8'd8  , 7'd91 , 2'd3, 2'd0};   //note: 7D
    assign memory[311] = {7'd69 , 8'd8  , 7'd91 , 2'd3, 2'd0};   //note: 7F
    assign memory[312] = {7'd66 , 8'd8  , 7'd91 , 2'd3, 2'd0};   //note: 7D
    assign memory[313] = {7'd69 , 8'd12 , 7'd92 , 2'd3, 2'd0};   //note: 7F
    assign memory[314] = {7'd66 , 8'd12 , 7'd92 , 2'd3, 2'd0};   //note: 7D
    assign memory[315] = {7'd69 , 8'd12 , 7'd94 , 2'd3, 2'd0};   //note: 7F
    assign memory[316] = {7'd66 , 8'd12 , 7'd92 , 2'd3, 2'd0};   //note: 7D
    assign memory[317] = {7'd69 , 8'd16 , 7'd92 , 2'd3, 2'd0};   //note: 7F
    assign memory[318] = {7'd66 , 8'd16 , 7'd92 , 2'd3, 2'd0};   //note: 7D
    assign memory[319] = {7'd69 , 8'd16 , 7'd94 , 2'd3, 2'd0};   //note: 7F
    assign memory[320] = {7'd66 , 8'd16 , 7'd94 , 2'd3, 2'd0};   //note: 7D
    assign memory[321] = {7'd69 , 8'd20 , 7'd94 , 2'd3, 2'd0};   //note: 7F
    assign memory[322] = {7'd66 , 8'd20 , 7'd94 , 2'd3, 2'd0};   //note: 7D
    assign memory[323] = {7'd69 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 7F
    assign memory[324] = {7'd66 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 7D
    assign memory[325] = {7'd69 , 8'd24 , 7'd94 , 2'd3, 2'd0};   //note: 7F
    assign memory[326] = {7'd66 , 8'd16 , 7'd94 , 2'd3, 2'd0};   //note: 7D
    assign memory[327] = {7'd69 , 8'd32 , 7'd94 , 2'd3, 2'd0};   //note: 7F
    assign memory[328] = {7'd66 , 8'd32 , 7'd94 , 2'd3, 2'd0};   //note: 7D
    assign memory[329] = {7'd69 , 8'd32 , 7'd94 , 2'd3, 2'd0};   //note: 7F
    assign memory[330] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[331] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[332] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[333] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[334] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[335] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[336] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[337] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[338] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[339] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[340] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[341] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[342] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[343] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[344] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[345] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[346] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[347] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[348] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[349] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[350] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[351] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[352] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[353] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[354] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[355] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[356] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[357] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[358] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[359] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[360] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[361] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[362] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[363] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[364] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[365] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[366] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[367] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[368] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[369] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[370] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[371] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[372] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[373] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[374] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[375] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[376] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[377] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[378] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[379] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[380] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[381] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[382] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[383] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[384] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[385] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[386] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[387] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[388] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[389] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[390] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[391] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[392] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[393] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[394] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[395] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[396] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[397] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[398] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[399] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[400] = {7'd0  , 8'd54 , 7'd0  , 2'd0, 2'd0};
    assign memory[401] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s1+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s1+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+79 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+80 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+81 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+82 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+83 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+84 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+85 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+86 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+87 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+88 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+89 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+90 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+91 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+92 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+93 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+94 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+95 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+96 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+97 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+98 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+99 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+100] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+101] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+102] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+103] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+104] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+105] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+106] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+107] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+108] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+109] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+110] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+111] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+112] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+113] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+114] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+115] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+116] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+117] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+118] = {7'd0  , 8'd118, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+119] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s2+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s2+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+2  ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+3  ] = {7'd40 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 5C
    assign memory[s2+4  ] = {7'd40 , 8'd129, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+5  ] = {7'd36 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+6  ] = {7'd36 , 8'd129, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+7  ] = {7'd36 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+8  ] = {7'd36 , 8'd129, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+9  ] = {7'd35 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4G
    assign memory[s2+10 ] = {7'd35 , 8'd129, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+12 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+13 ] = {7'd33 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+14 ] = {7'd33 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+15 ] = {7'd33 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+16 ] = {7'd33 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+17 ] = {7'd31 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+18 ] = {7'd31 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+19 ] = {7'd31 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+20 ] = {7'd31 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+21 ] = {7'd33 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+22 ] = {7'd33 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+23 ] = {7'd33 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+24 ] = {7'd33 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+25 ] = {7'd31 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+26 ] = {7'd31 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+27 ] = {7'd31 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+28 ] = {7'd31 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+29 ] = {7'd36 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+30 ] = {7'd36 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+31 ] = {7'd36 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+32 ] = {7'd36 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+33 ] = {7'd36 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+34 ] = {7'd36 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+35 ] = {7'd35 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4G
    assign memory[s2+36 ] = {7'd35 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+37 ] = {7'd36 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+38 ] = {7'd36 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+39 ] = {7'd36 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+40 ] = {7'd36 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+41 ] = {7'd36 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+42 ] = {7'd36 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+43 ] = {7'd35 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4G
    assign memory[s2+44 ] = {7'd35 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+45 ] = {7'd40 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 5C
    assign memory[s2+46 ] = {7'd40 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+47 ] = {7'd41 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s2+48 ] = {7'd41 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+49 ] = {7'd36 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+50 ] = {7'd36 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+52 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+53 ] = {7'd40 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 5C
    assign memory[s2+54 ] = {7'd40 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+55 ] = {7'd41 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s2+56 ] = {7'd41 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+57 ] = {7'd40 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 5C
    assign memory[s2+58 ] = {7'd40 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+59 ] = {7'd38 , 8'd192, 7'd95 , 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s2+60 ] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+61 ] = {7'd40 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 5C
    assign memory[s2+62 ] = {7'd40 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+63 ] = {7'd40 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 5C
    assign memory[s2+64 ] = {7'd36 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+65 ] = {7'd36 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+66 ] = {7'd36 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+67 ] = {7'd36 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+68 ] = {7'd36 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+69 ] = {7'd36 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+70 ] = {7'd35 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G
    assign memory[s2+71 ] = {7'd35 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+72 ] = {7'd35 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G
    assign memory[s2+73 ] = {7'd40 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 5C
    assign memory[s2+74 ] = {7'd40 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+75 ] = {7'd40 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 5C
    assign memory[s2+76 ] = {7'd36 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+77 ] = {7'd36 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+78 ] = {7'd36 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+79 ] = {7'd36 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+80 ] = {7'd36 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+81 ] = {7'd36 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+82 ] = {7'd35 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G
    assign memory[s2+83 ] = {7'd35 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+84 ] = {7'd35 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G
    assign memory[s2+85 ] = {7'd40 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 5C
    assign memory[s2+86 ] = {7'd40 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+87 ] = {7'd40 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 5C
    assign memory[s2+88 ] = {7'd36 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+89 ] = {7'd36 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+90 ] = {7'd36 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+91 ] = {7'd36 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+92 ] = {7'd36 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+93 ] = {7'd36 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+94 ] = {7'd35 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G
    assign memory[s2+95 ] = {7'd35 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+96 ] = {7'd35 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G
    assign memory[s2+97 ] = {7'd40 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 5C
    assign memory[s2+98 ] = {7'd40 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+99 ] = {7'd40 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 5C
    assign memory[s2+100] = {7'd36 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+101] = {7'd36 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+102] = {7'd36 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+103] = {7'd36 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+104] = {7'd36 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+105] = {7'd36 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+106] = {7'd35 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4G
    assign memory[s2+107] = {7'd35 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s2+108] = {7'd40 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 5C
    assign memory[s2+109] = {7'd40 , 8'd33 , 7'd72 , 2'd0, 2'd0};
    assign memory[s2+110] = {7'd40 , 8'd96 , 7'd72 , 2'd0, 2'd0};   //note: 5C
    assign memory[s2+111] = {7'd36 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+112] = {7'd36 , 8'd33 , 7'd72 , 2'd0, 2'd0};
    assign memory[s2+113] = {7'd36 , 8'd96 , 7'd72 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+114] = {7'd36 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+115] = {7'd36 , 8'd33 , 7'd72 , 2'd0, 2'd0};
    assign memory[s2+116] = {7'd36 , 8'd96 , 7'd72 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+117] = {7'd35 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4G
    assign memory[s2+118] = {7'd35 , 8'd255, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+119] = {7'd35 , 8'd66 , 7'd72 , 2'd0, 2'd0};
    assign memory[s2+120] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+121] = {7'd0  , 8'd1  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+122] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+123] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+124] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s3+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s3+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+13 ] = {7'd0  , 8'd112, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+14 ] = {7'd32 , 8'd184, 7'd79 , 2'd0, 2'd0};   //note: 4E
    assign memory[s3+15 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+16 ] = {7'd31 , 8'd184, 7'd79 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+17 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+18 ] = {7'd34 , 8'd184, 7'd79 , 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s3+19 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+20 ] = {7'd31 , 8'd184, 7'd79 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+21 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+22 ] = {7'd32 , 8'd184, 7'd79 , 2'd0, 2'd0};   //note: 4E
    assign memory[s3+23 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+24 ] = {7'd31 , 8'd184, 7'd79 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+25 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+26 ] = {7'd34 , 8'd184, 7'd79 , 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s3+27 ] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+28 ] = {7'd31 , 8'd92 , 7'd79 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+54 ] = {7'd0  , 8'd57 , 7'd0  , 2'd0, 2'd0};
    assign memory[s3+55 ] = {7'd40 , 8'd192, 7'd101, 2'd0, 2'd0};   //note: 5C
    assign memory[s3+56 ] = {7'd36 , 8'd192, 7'd98 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s3+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+59 ] = {7'd0  , 8'd66 , 7'd0  , 2'd0, 2'd0};
    assign memory[s3+60 ] = {7'd33 , 8'd48 , 7'd88 , 2'd0, 2'd0};   //note: 4F
    assign memory[s3+61 ] = {7'd35 , 8'd48 , 7'd88 , 2'd0, 2'd0};   //note: 4G
    assign memory[s3+62 ] = {7'd36 , 8'd48 , 7'd88 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s3+63 ] = {7'd38 , 8'd48 , 7'd88 , 2'd0, 2'd0};   //note: 4A#Bb
    assign memory[s3+64 ] = {7'd39 , 8'd48 , 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+65 ] = {7'd39 , 8'd48 , 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+66 ] = {7'd41 , 8'd48 , 7'd88 , 2'd0, 2'd0};   //note: 5C#Db
    assign memory[s3+67 ] = {7'd43 , 8'd48 , 7'd88 , 2'd0, 2'd0};   //note: 5D#Eb
    assign memory[s3+68 ] = {7'd44 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 5E
    assign memory[s3+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+79 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+80 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+81 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+82 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+83 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+84 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+85 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+86 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+87 ] = {7'd0  , 8'd114, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+88 ] = {7'd51 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 5B
    assign memory[s3+89 ] = {7'd51 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 5B
    assign memory[s3+90 ] = {7'd51 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 5B
    assign memory[s3+91 ] = {7'd51 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 5B
    assign memory[s3+92 ] = {7'd51 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 5B
    assign memory[s3+93 ] = {7'd51 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 5B
    assign memory[s3+94 ] = {7'd51 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 5B
    assign memory[s3+95 ] = {7'd51 , 8'd255, 7'd88 , 2'd0, 2'd0};   //note: 5B
    assign memory[s3+96 ] = {7'd51 , 8'd225, 7'd88 , 2'd0, 2'd0};
    assign memory[s3+97 ] = {7'd0  , 8'd2  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+98 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+99 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+100] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song


endmodule							
