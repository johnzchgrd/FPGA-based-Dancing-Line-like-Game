`timescale 1ns / 1ps

module hint_songsel_rom(
   input valid,
   input [8:0]x,
   input [4:0]y,
   output reg songsel_type
    );
    wire memhint[8578:0];
    always @(*)begin
        if(valid)begin
            songsel_type = memhint[x+y*373];
        end else begin
            songsel_type = 1'b0;
        end
    end
    
    assign memhint[0   ] = 1'd0;
    assign memhint[1   ] = 1'd0;
    assign memhint[2   ] = 1'd0;
    assign memhint[3   ] = 1'd0;
    assign memhint[4   ] = 1'd1;
    assign memhint[5   ] = 1'd1;
    assign memhint[6   ] = 1'd1;
    assign memhint[7   ] = 1'd1;
    assign memhint[8   ] = 1'd1;
    assign memhint[9   ] = 1'd0;
    assign memhint[10  ] = 1'd0;
    assign memhint[11  ] = 1'd0;
    assign memhint[12  ] = 1'd0;
    assign memhint[13  ] = 1'd0;
    assign memhint[14  ] = 1'd0;
    assign memhint[15  ] = 1'd0;
    assign memhint[16  ] = 1'd0;
    assign memhint[17  ] = 1'd0;
    assign memhint[18  ] = 1'd1;
    assign memhint[19  ] = 1'd1;
    assign memhint[20  ] = 1'd1;
    assign memhint[21  ] = 1'd1;
    assign memhint[22  ] = 1'd1;
    assign memhint[23  ] = 1'd1;
    assign memhint[24  ] = 1'd1;
    assign memhint[25  ] = 1'd1;
    assign memhint[26  ] = 1'd1;
    assign memhint[27  ] = 1'd1;
    assign memhint[28  ] = 1'd1;
    assign memhint[29  ] = 1'd1;
    assign memhint[30  ] = 1'd1;
    assign memhint[31  ] = 1'd0;
    assign memhint[32  ] = 1'd0;
    assign memhint[33  ] = 1'd0;
    assign memhint[34  ] = 1'd0;
    assign memhint[35  ] = 1'd1;
    assign memhint[36  ] = 1'd1;
    assign memhint[37  ] = 1'd0;
    assign memhint[38  ] = 1'd0;
    assign memhint[39  ] = 1'd0;
    assign memhint[40  ] = 1'd0;
    assign memhint[41  ] = 1'd0;
    assign memhint[42  ] = 1'd0;
    assign memhint[43  ] = 1'd0;
    assign memhint[44  ] = 1'd0;
    assign memhint[45  ] = 1'd0;
    assign memhint[46  ] = 1'd0;
    assign memhint[47  ] = 1'd0;
    assign memhint[48  ] = 1'd0;
    assign memhint[49  ] = 1'd0;
    assign memhint[50  ] = 1'd1;
    assign memhint[51  ] = 1'd1;
    assign memhint[52  ] = 1'd1;
    assign memhint[53  ] = 1'd1;
    assign memhint[54  ] = 1'd1;
    assign memhint[55  ] = 1'd1;
    assign memhint[56  ] = 1'd1;
    assign memhint[57  ] = 1'd1;
    assign memhint[58  ] = 1'd1;
    assign memhint[59  ] = 1'd1;
    assign memhint[60  ] = 1'd1;
    assign memhint[61  ] = 1'd1;
    assign memhint[62  ] = 1'd1;
    assign memhint[63  ] = 1'd0;
    assign memhint[64  ] = 1'd0;
    assign memhint[65  ] = 1'd0;
    assign memhint[66  ] = 1'd0;
    assign memhint[67  ] = 1'd0;
    assign memhint[68  ] = 1'd0;
    assign memhint[69  ] = 1'd0;
    assign memhint[70  ] = 1'd0;
    assign memhint[71  ] = 1'd0;
    assign memhint[72  ] = 1'd0;
    assign memhint[73  ] = 1'd0;
    assign memhint[74  ] = 1'd1;
    assign memhint[75  ] = 1'd1;
    assign memhint[76  ] = 1'd1;
    assign memhint[77  ] = 1'd1;
    assign memhint[78  ] = 1'd1;
    assign memhint[79  ] = 1'd1;
    assign memhint[80  ] = 1'd1;
    assign memhint[81  ] = 1'd1;
    assign memhint[82  ] = 1'd0;
    assign memhint[83  ] = 1'd0;
    assign memhint[84  ] = 1'd0;
    assign memhint[85  ] = 1'd0;
    assign memhint[86  ] = 1'd0;
    assign memhint[87  ] = 1'd0;
    assign memhint[88  ] = 1'd0;
    assign memhint[89  ] = 1'd0;
    assign memhint[90  ] = 1'd1;
    assign memhint[91  ] = 1'd1;
    assign memhint[92  ] = 1'd1;
    assign memhint[93  ] = 1'd1;
    assign memhint[94  ] = 1'd1;
    assign memhint[95  ] = 1'd1;
    assign memhint[96  ] = 1'd1;
    assign memhint[97  ] = 1'd1;
    assign memhint[98  ] = 1'd1;
    assign memhint[99  ] = 1'd1;
    assign memhint[100 ] = 1'd1;
    assign memhint[101 ] = 1'd1;
    assign memhint[102 ] = 1'd0;
    assign memhint[103 ] = 1'd0;
    assign memhint[104 ] = 1'd0;
    assign memhint[105 ] = 1'd0;
    assign memhint[106 ] = 1'd0;
    assign memhint[107 ] = 1'd0;
    assign memhint[108 ] = 1'd0;
    assign memhint[109 ] = 1'd0;
    assign memhint[110 ] = 1'd0;
    assign memhint[111 ] = 1'd0;
    assign memhint[112 ] = 1'd0;
    assign memhint[113 ] = 1'd0;
    assign memhint[114 ] = 1'd0;
    assign memhint[115 ] = 1'd0;
    assign memhint[116 ] = 1'd0;
    assign memhint[117 ] = 1'd0;
    assign memhint[118 ] = 1'd0;
    assign memhint[119 ] = 1'd0;
    assign memhint[120 ] = 1'd0;
    assign memhint[121 ] = 1'd0;
    assign memhint[122 ] = 1'd0;
    assign memhint[123 ] = 1'd1;
    assign memhint[124 ] = 1'd0;
    assign memhint[125 ] = 1'd0;
    assign memhint[126 ] = 1'd0;
    assign memhint[127 ] = 1'd0;
    assign memhint[128 ] = 1'd0;
    assign memhint[129 ] = 1'd0;
    assign memhint[130 ] = 1'd0;
    assign memhint[131 ] = 1'd0;
    assign memhint[132 ] = 1'd0;
    assign memhint[133 ] = 1'd0;
    assign memhint[134 ] = 1'd0;
    assign memhint[135 ] = 1'd0;
    assign memhint[136 ] = 1'd0;
    assign memhint[137 ] = 1'd0;
    assign memhint[138 ] = 1'd0;
    assign memhint[139 ] = 1'd0;
    assign memhint[140 ] = 1'd0;
    assign memhint[141 ] = 1'd0;
    assign memhint[142 ] = 1'd0;
    assign memhint[143 ] = 1'd0;
    assign memhint[144 ] = 1'd0;
    assign memhint[145 ] = 1'd0;
    assign memhint[146 ] = 1'd0;
    assign memhint[147 ] = 1'd0;
    assign memhint[148 ] = 1'd0;
    assign memhint[149 ] = 1'd1;
    assign memhint[150 ] = 1'd1;
    assign memhint[151 ] = 1'd1;
    assign memhint[152 ] = 1'd1;
    assign memhint[153 ] = 1'd1;
    assign memhint[154 ] = 1'd0;
    assign memhint[155 ] = 1'd0;
    assign memhint[156 ] = 1'd0;
    assign memhint[157 ] = 1'd0;
    assign memhint[158 ] = 1'd0;
    assign memhint[159 ] = 1'd0;
    assign memhint[160 ] = 1'd0;
    assign memhint[161 ] = 1'd0;
    assign memhint[162 ] = 1'd0;
    assign memhint[163 ] = 1'd0;
    assign memhint[164 ] = 1'd0;
    assign memhint[165 ] = 1'd0;
    assign memhint[166 ] = 1'd0;
    assign memhint[167 ] = 1'd0;
    assign memhint[168 ] = 1'd0;
    assign memhint[169 ] = 1'd0;
    assign memhint[170 ] = 1'd1;
    assign memhint[171 ] = 1'd1;
    assign memhint[172 ] = 1'd1;
    assign memhint[173 ] = 1'd1;
    assign memhint[174 ] = 1'd1;
    assign memhint[175 ] = 1'd1;
    assign memhint[176 ] = 1'd1;
    assign memhint[177 ] = 1'd1;
    assign memhint[178 ] = 1'd0;
    assign memhint[179 ] = 1'd0;
    assign memhint[180 ] = 1'd0;
    assign memhint[181 ] = 1'd0;
    assign memhint[182 ] = 1'd0;
    assign memhint[183 ] = 1'd0;
    assign memhint[184 ] = 1'd0;
    assign memhint[185 ] = 1'd0;
    assign memhint[186 ] = 1'd0;
    assign memhint[187 ] = 1'd0;
    assign memhint[188 ] = 1'd0;
    assign memhint[189 ] = 1'd0;
    assign memhint[190 ] = 1'd0;
    assign memhint[191 ] = 1'd1;
    assign memhint[192 ] = 1'd0;
    assign memhint[193 ] = 1'd0;
    assign memhint[194 ] = 1'd0;
    assign memhint[195 ] = 1'd0;
    assign memhint[196 ] = 1'd0;
    assign memhint[197 ] = 1'd0;
    assign memhint[198 ] = 1'd0;
    assign memhint[199 ] = 1'd0;
    assign memhint[200 ] = 1'd0;
    assign memhint[201 ] = 1'd0;
    assign memhint[202 ] = 1'd0;
    assign memhint[203 ] = 1'd0;
    assign memhint[204 ] = 1'd0;
    assign memhint[205 ] = 1'd0;
    assign memhint[206 ] = 1'd0;
    assign memhint[207 ] = 1'd1;
    assign memhint[208 ] = 1'd1;
    assign memhint[209 ] = 1'd0;
    assign memhint[210 ] = 1'd0;
    assign memhint[211 ] = 1'd0;
    assign memhint[212 ] = 1'd0;
    assign memhint[213 ] = 1'd0;
    assign memhint[214 ] = 1'd0;
    assign memhint[215 ] = 1'd0;
    assign memhint[216 ] = 1'd0;
    assign memhint[217 ] = 1'd0;
    assign memhint[218 ] = 1'd0;
    assign memhint[219 ] = 1'd0;
    assign memhint[220 ] = 1'd0;
    assign memhint[221 ] = 1'd0;
    assign memhint[222 ] = 1'd0;
    assign memhint[223 ] = 1'd1;
    assign memhint[224 ] = 1'd1;
    assign memhint[225 ] = 1'd1;
    assign memhint[226 ] = 1'd1;
    assign memhint[227 ] = 1'd1;
    assign memhint[228 ] = 1'd1;
    assign memhint[229 ] = 1'd1;
    assign memhint[230 ] = 1'd0;
    assign memhint[231 ] = 1'd0;
    assign memhint[232 ] = 1'd0;
    assign memhint[233 ] = 1'd0;
    assign memhint[234 ] = 1'd0;
    assign memhint[235 ] = 1'd0;
    assign memhint[236 ] = 1'd0;
    assign memhint[237 ] = 1'd0;
    assign memhint[238 ] = 1'd0;
    assign memhint[239 ] = 1'd0;
    assign memhint[240 ] = 1'd0;
    assign memhint[241 ] = 1'd0;
    assign memhint[242 ] = 1'd0;
    assign memhint[243 ] = 1'd0;
    assign memhint[244 ] = 1'd0;
    assign memhint[245 ] = 1'd0;
    assign memhint[246 ] = 1'd0;
    assign memhint[247 ] = 1'd0;
    assign memhint[248 ] = 1'd0;
    assign memhint[249 ] = 1'd1;
    assign memhint[250 ] = 1'd1;
    assign memhint[251 ] = 1'd1;
    assign memhint[252 ] = 1'd1;
    assign memhint[253 ] = 1'd1;
    assign memhint[254 ] = 1'd1;
    assign memhint[255 ] = 1'd1;
    assign memhint[256 ] = 1'd1;
    assign memhint[257 ] = 1'd1;
    assign memhint[258 ] = 1'd1;
    assign memhint[259 ] = 1'd1;
    assign memhint[260 ] = 1'd1;
    assign memhint[261 ] = 1'd0;
    assign memhint[262 ] = 1'd0;
    assign memhint[263 ] = 1'd0;
    assign memhint[264 ] = 1'd0;
    assign memhint[265 ] = 1'd0;
    assign memhint[266 ] = 1'd0;
    assign memhint[267 ] = 1'd0;
    assign memhint[268 ] = 1'd0;
    assign memhint[269 ] = 1'd0;
    assign memhint[270 ] = 1'd0;
    assign memhint[271 ] = 1'd0;
    assign memhint[272 ] = 1'd1;
    assign memhint[273 ] = 1'd1;
    assign memhint[274 ] = 1'd1;
    assign memhint[275 ] = 1'd1;
    assign memhint[276 ] = 1'd1;
    assign memhint[277 ] = 1'd1;
    assign memhint[278 ] = 1'd1;
    assign memhint[279 ] = 1'd1;
    assign memhint[280 ] = 1'd0;
    assign memhint[281 ] = 1'd0;
    assign memhint[282 ] = 1'd0;
    assign memhint[283 ] = 1'd0;
    assign memhint[284 ] = 1'd0;
    assign memhint[285 ] = 1'd0;
    assign memhint[286 ] = 1'd0;
    assign memhint[287 ] = 1'd0;
    assign memhint[288 ] = 1'd0;
    assign memhint[289 ] = 1'd0;
    assign memhint[290 ] = 1'd0;
    assign memhint[291 ] = 1'd0;
    assign memhint[292 ] = 1'd0;
    assign memhint[293 ] = 1'd0;
    assign memhint[294 ] = 1'd0;
    assign memhint[295 ] = 1'd0;
    assign memhint[296 ] = 1'd0;
    assign memhint[297 ] = 1'd0;
    assign memhint[298 ] = 1'd0;
    assign memhint[299 ] = 1'd0;
    assign memhint[300 ] = 1'd0;
    assign memhint[301 ] = 1'd0;
    assign memhint[302 ] = 1'd1;
    assign memhint[303 ] = 1'd1;
    assign memhint[304 ] = 1'd1;
    assign memhint[305 ] = 1'd1;
    assign memhint[306 ] = 1'd1;
    assign memhint[307 ] = 1'd1;
    assign memhint[308 ] = 1'd1;
    assign memhint[309 ] = 1'd1;
    assign memhint[310 ] = 1'd1;
    assign memhint[311 ] = 1'd1;
    assign memhint[312 ] = 1'd0;
    assign memhint[313 ] = 1'd0;
    assign memhint[314 ] = 1'd0;
    assign memhint[315 ] = 1'd0;
    assign memhint[316 ] = 1'd0;
    assign memhint[317 ] = 1'd0;
    assign memhint[318 ] = 1'd0;
    assign memhint[319 ] = 1'd0;
    assign memhint[320 ] = 1'd0;
    assign memhint[321 ] = 1'd1;
    assign memhint[322 ] = 1'd1;
    assign memhint[323 ] = 1'd0;
    assign memhint[324 ] = 1'd0;
    assign memhint[325 ] = 1'd0;
    assign memhint[326 ] = 1'd0;
    assign memhint[327 ] = 1'd0;
    assign memhint[328 ] = 1'd0;
    assign memhint[329 ] = 1'd0;
    assign memhint[330 ] = 1'd0;
    assign memhint[331 ] = 1'd0;
    assign memhint[332 ] = 1'd0;
    assign memhint[333 ] = 1'd0;
    assign memhint[334 ] = 1'd0;
    assign memhint[335 ] = 1'd0;
    assign memhint[336 ] = 1'd0;
    assign memhint[337 ] = 1'd0;
    assign memhint[338 ] = 1'd0;
    assign memhint[339 ] = 1'd0;
    assign memhint[340 ] = 1'd0;
    assign memhint[341 ] = 1'd0;
    assign memhint[342 ] = 1'd0;
    assign memhint[343 ] = 1'd0;
    assign memhint[344 ] = 1'd1;
    assign memhint[345 ] = 1'd0;
    assign memhint[346 ] = 1'd0;
    assign memhint[347 ] = 1'd0;
    assign memhint[348 ] = 1'd0;
    assign memhint[349 ] = 1'd0;
    assign memhint[350 ] = 1'd0;
    assign memhint[351 ] = 1'd0;
    assign memhint[352 ] = 1'd0;
    assign memhint[353 ] = 1'd0;
    assign memhint[354 ] = 1'd0;
    assign memhint[355 ] = 1'd0;
    assign memhint[356 ] = 1'd0;
    assign memhint[357 ] = 1'd1;
    assign memhint[358 ] = 1'd1;
    assign memhint[359 ] = 1'd0;
    assign memhint[360 ] = 1'd0;
    assign memhint[361 ] = 1'd0;
    assign memhint[362 ] = 1'd0;
    assign memhint[363 ] = 1'd0;
    assign memhint[364 ] = 1'd0;
    assign memhint[365 ] = 1'd0;
    assign memhint[366 ] = 1'd0;
    assign memhint[367 ] = 1'd0;
    assign memhint[368 ] = 1'd0;
    assign memhint[369 ] = 1'd0;
    assign memhint[370 ] = 1'd0;
    assign memhint[371 ] = 1'd1;
    assign memhint[372 ] = 1'd1;
    assign memhint[373 ] = 1'd0;
    assign memhint[374 ] = 1'd0;
    assign memhint[375 ] = 1'd0;
    assign memhint[376 ] = 1'd1;
    assign memhint[377 ] = 1'd1;
    assign memhint[378 ] = 1'd1;
    assign memhint[379 ] = 1'd1;
    assign memhint[380 ] = 1'd1;
    assign memhint[381 ] = 1'd1;
    assign memhint[382 ] = 1'd1;
    assign memhint[383 ] = 1'd1;
    assign memhint[384 ] = 1'd0;
    assign memhint[385 ] = 1'd0;
    assign memhint[386 ] = 1'd0;
    assign memhint[387 ] = 1'd0;
    assign memhint[388 ] = 1'd0;
    assign memhint[389 ] = 1'd0;
    assign memhint[390 ] = 1'd0;
    assign memhint[391 ] = 1'd1;
    assign memhint[392 ] = 1'd1;
    assign memhint[393 ] = 1'd1;
    assign memhint[394 ] = 1'd1;
    assign memhint[395 ] = 1'd1;
    assign memhint[396 ] = 1'd1;
    assign memhint[397 ] = 1'd1;
    assign memhint[398 ] = 1'd1;
    assign memhint[399 ] = 1'd1;
    assign memhint[400 ] = 1'd1;
    assign memhint[401 ] = 1'd1;
    assign memhint[402 ] = 1'd1;
    assign memhint[403 ] = 1'd1;
    assign memhint[404 ] = 1'd0;
    assign memhint[405 ] = 1'd0;
    assign memhint[406 ] = 1'd0;
    assign memhint[407 ] = 1'd0;
    assign memhint[408 ] = 1'd1;
    assign memhint[409 ] = 1'd1;
    assign memhint[410 ] = 1'd0;
    assign memhint[411 ] = 1'd0;
    assign memhint[412 ] = 1'd0;
    assign memhint[413 ] = 1'd0;
    assign memhint[414 ] = 1'd0;
    assign memhint[415 ] = 1'd0;
    assign memhint[416 ] = 1'd0;
    assign memhint[417 ] = 1'd0;
    assign memhint[418 ] = 1'd0;
    assign memhint[419 ] = 1'd0;
    assign memhint[420 ] = 1'd0;
    assign memhint[421 ] = 1'd0;
    assign memhint[422 ] = 1'd0;
    assign memhint[423 ] = 1'd1;
    assign memhint[424 ] = 1'd1;
    assign memhint[425 ] = 1'd1;
    assign memhint[426 ] = 1'd1;
    assign memhint[427 ] = 1'd1;
    assign memhint[428 ] = 1'd1;
    assign memhint[429 ] = 1'd1;
    assign memhint[430 ] = 1'd1;
    assign memhint[431 ] = 1'd1;
    assign memhint[432 ] = 1'd1;
    assign memhint[433 ] = 1'd1;
    assign memhint[434 ] = 1'd1;
    assign memhint[435 ] = 1'd1;
    assign memhint[436 ] = 1'd0;
    assign memhint[437 ] = 1'd0;
    assign memhint[438 ] = 1'd0;
    assign memhint[439 ] = 1'd0;
    assign memhint[440 ] = 1'd0;
    assign memhint[441 ] = 1'd0;
    assign memhint[442 ] = 1'd0;
    assign memhint[443 ] = 1'd0;
    assign memhint[444 ] = 1'd0;
    assign memhint[445 ] = 1'd1;
    assign memhint[446 ] = 1'd1;
    assign memhint[447 ] = 1'd1;
    assign memhint[448 ] = 1'd1;
    assign memhint[449 ] = 1'd1;
    assign memhint[450 ] = 1'd1;
    assign memhint[451 ] = 1'd1;
    assign memhint[452 ] = 1'd1;
    assign memhint[453 ] = 1'd1;
    assign memhint[454 ] = 1'd1;
    assign memhint[455 ] = 1'd1;
    assign memhint[456 ] = 1'd1;
    assign memhint[457 ] = 1'd0;
    assign memhint[458 ] = 1'd0;
    assign memhint[459 ] = 1'd0;
    assign memhint[460 ] = 1'd0;
    assign memhint[461 ] = 1'd0;
    assign memhint[462 ] = 1'd0;
    assign memhint[463 ] = 1'd1;
    assign memhint[464 ] = 1'd1;
    assign memhint[465 ] = 1'd1;
    assign memhint[466 ] = 1'd1;
    assign memhint[467 ] = 1'd1;
    assign memhint[468 ] = 1'd1;
    assign memhint[469 ] = 1'd1;
    assign memhint[470 ] = 1'd1;
    assign memhint[471 ] = 1'd1;
    assign memhint[472 ] = 1'd1;
    assign memhint[473 ] = 1'd1;
    assign memhint[474 ] = 1'd1;
    assign memhint[475 ] = 1'd0;
    assign memhint[476 ] = 1'd0;
    assign memhint[477 ] = 1'd0;
    assign memhint[478 ] = 1'd0;
    assign memhint[479 ] = 1'd0;
    assign memhint[480 ] = 1'd0;
    assign memhint[481 ] = 1'd0;
    assign memhint[482 ] = 1'd0;
    assign memhint[483 ] = 1'd0;
    assign memhint[484 ] = 1'd0;
    assign memhint[485 ] = 1'd0;
    assign memhint[486 ] = 1'd0;
    assign memhint[487 ] = 1'd0;
    assign memhint[488 ] = 1'd0;
    assign memhint[489 ] = 1'd0;
    assign memhint[490 ] = 1'd0;
    assign memhint[491 ] = 1'd0;
    assign memhint[492 ] = 1'd0;
    assign memhint[493 ] = 1'd0;
    assign memhint[494 ] = 1'd0;
    assign memhint[495 ] = 1'd1;
    assign memhint[496 ] = 1'd1;
    assign memhint[497 ] = 1'd1;
    assign memhint[498 ] = 1'd0;
    assign memhint[499 ] = 1'd0;
    assign memhint[500 ] = 1'd0;
    assign memhint[501 ] = 1'd0;
    assign memhint[502 ] = 1'd0;
    assign memhint[503 ] = 1'd0;
    assign memhint[504 ] = 1'd0;
    assign memhint[505 ] = 1'd0;
    assign memhint[506 ] = 1'd0;
    assign memhint[507 ] = 1'd0;
    assign memhint[508 ] = 1'd0;
    assign memhint[509 ] = 1'd0;
    assign memhint[510 ] = 1'd0;
    assign memhint[511 ] = 1'd0;
    assign memhint[512 ] = 1'd0;
    assign memhint[513 ] = 1'd0;
    assign memhint[514 ] = 1'd0;
    assign memhint[515 ] = 1'd0;
    assign memhint[516 ] = 1'd0;
    assign memhint[517 ] = 1'd0;
    assign memhint[518 ] = 1'd0;
    assign memhint[519 ] = 1'd0;
    assign memhint[520 ] = 1'd0;
    assign memhint[521 ] = 1'd1;
    assign memhint[522 ] = 1'd1;
    assign memhint[523 ] = 1'd1;
    assign memhint[524 ] = 1'd1;
    assign memhint[525 ] = 1'd1;
    assign memhint[526 ] = 1'd1;
    assign memhint[527 ] = 1'd1;
    assign memhint[528 ] = 1'd1;
    assign memhint[529 ] = 1'd0;
    assign memhint[530 ] = 1'd0;
    assign memhint[531 ] = 1'd0;
    assign memhint[532 ] = 1'd0;
    assign memhint[533 ] = 1'd0;
    assign memhint[534 ] = 1'd0;
    assign memhint[535 ] = 1'd0;
    assign memhint[536 ] = 1'd0;
    assign memhint[537 ] = 1'd0;
    assign memhint[538 ] = 1'd0;
    assign memhint[539 ] = 1'd0;
    assign memhint[540 ] = 1'd0;
    assign memhint[541 ] = 1'd1;
    assign memhint[542 ] = 1'd1;
    assign memhint[543 ] = 1'd1;
    assign memhint[544 ] = 1'd1;
    assign memhint[545 ] = 1'd1;
    assign memhint[546 ] = 1'd1;
    assign memhint[547 ] = 1'd1;
    assign memhint[548 ] = 1'd1;
    assign memhint[549 ] = 1'd1;
    assign memhint[550 ] = 1'd1;
    assign memhint[551 ] = 1'd1;
    assign memhint[552 ] = 1'd1;
    assign memhint[553 ] = 1'd0;
    assign memhint[554 ] = 1'd0;
    assign memhint[555 ] = 1'd0;
    assign memhint[556 ] = 1'd0;
    assign memhint[557 ] = 1'd0;
    assign memhint[558 ] = 1'd0;
    assign memhint[559 ] = 1'd0;
    assign memhint[560 ] = 1'd0;
    assign memhint[561 ] = 1'd0;
    assign memhint[562 ] = 1'd0;
    assign memhint[563 ] = 1'd0;
    assign memhint[564 ] = 1'd1;
    assign memhint[565 ] = 1'd1;
    assign memhint[566 ] = 1'd0;
    assign memhint[567 ] = 1'd0;
    assign memhint[568 ] = 1'd0;
    assign memhint[569 ] = 1'd0;
    assign memhint[570 ] = 1'd0;
    assign memhint[571 ] = 1'd0;
    assign memhint[572 ] = 1'd0;
    assign memhint[573 ] = 1'd0;
    assign memhint[574 ] = 1'd0;
    assign memhint[575 ] = 1'd0;
    assign memhint[576 ] = 1'd0;
    assign memhint[577 ] = 1'd0;
    assign memhint[578 ] = 1'd0;
    assign memhint[579 ] = 1'd0;
    assign memhint[580 ] = 1'd1;
    assign memhint[581 ] = 1'd1;
    assign memhint[582 ] = 1'd0;
    assign memhint[583 ] = 1'd0;
    assign memhint[584 ] = 1'd0;
    assign memhint[585 ] = 1'd0;
    assign memhint[586 ] = 1'd0;
    assign memhint[587 ] = 1'd0;
    assign memhint[588 ] = 1'd0;
    assign memhint[589 ] = 1'd0;
    assign memhint[590 ] = 1'd0;
    assign memhint[591 ] = 1'd0;
    assign memhint[592 ] = 1'd0;
    assign memhint[593 ] = 1'd1;
    assign memhint[594 ] = 1'd1;
    assign memhint[595 ] = 1'd1;
    assign memhint[596 ] = 1'd1;
    assign memhint[597 ] = 1'd1;
    assign memhint[598 ] = 1'd1;
    assign memhint[599 ] = 1'd1;
    assign memhint[600 ] = 1'd1;
    assign memhint[601 ] = 1'd1;
    assign memhint[602 ] = 1'd1;
    assign memhint[603 ] = 1'd1;
    assign memhint[604 ] = 1'd1;
    assign memhint[605 ] = 1'd1;
    assign memhint[606 ] = 1'd0;
    assign memhint[607 ] = 1'd0;
    assign memhint[608 ] = 1'd0;
    assign memhint[609 ] = 1'd0;
    assign memhint[610 ] = 1'd0;
    assign memhint[611 ] = 1'd0;
    assign memhint[612 ] = 1'd0;
    assign memhint[613 ] = 1'd0;
    assign memhint[614 ] = 1'd0;
    assign memhint[615 ] = 1'd0;
    assign memhint[616 ] = 1'd0;
    assign memhint[617 ] = 1'd0;
    assign memhint[618 ] = 1'd0;
    assign memhint[619 ] = 1'd0;
    assign memhint[620 ] = 1'd0;
    assign memhint[621 ] = 1'd0;
    assign memhint[622 ] = 1'd1;
    assign memhint[623 ] = 1'd1;
    assign memhint[624 ] = 1'd1;
    assign memhint[625 ] = 1'd1;
    assign memhint[626 ] = 1'd1;
    assign memhint[627 ] = 1'd1;
    assign memhint[628 ] = 1'd1;
    assign memhint[629 ] = 1'd1;
    assign memhint[630 ] = 1'd1;
    assign memhint[631 ] = 1'd1;
    assign memhint[632 ] = 1'd1;
    assign memhint[633 ] = 1'd1;
    assign memhint[634 ] = 1'd0;
    assign memhint[635 ] = 1'd0;
    assign memhint[636 ] = 1'd0;
    assign memhint[637 ] = 1'd0;
    assign memhint[638 ] = 1'd0;
    assign memhint[639 ] = 1'd0;
    assign memhint[640 ] = 1'd0;
    assign memhint[641 ] = 1'd0;
    assign memhint[642 ] = 1'd0;
    assign memhint[643 ] = 1'd1;
    assign memhint[644 ] = 1'd1;
    assign memhint[645 ] = 1'd1;
    assign memhint[646 ] = 1'd1;
    assign memhint[647 ] = 1'd1;
    assign memhint[648 ] = 1'd1;
    assign memhint[649 ] = 1'd1;
    assign memhint[650 ] = 1'd1;
    assign memhint[651 ] = 1'd1;
    assign memhint[652 ] = 1'd1;
    assign memhint[653 ] = 1'd1;
    assign memhint[654 ] = 1'd1;
    assign memhint[655 ] = 1'd0;
    assign memhint[656 ] = 1'd0;
    assign memhint[657 ] = 1'd0;
    assign memhint[658 ] = 1'd0;
    assign memhint[659 ] = 1'd0;
    assign memhint[660 ] = 1'd0;
    assign memhint[661 ] = 1'd0;
    assign memhint[662 ] = 1'd0;
    assign memhint[663 ] = 1'd0;
    assign memhint[664 ] = 1'd0;
    assign memhint[665 ] = 1'd0;
    assign memhint[666 ] = 1'd0;
    assign memhint[667 ] = 1'd0;
    assign memhint[668 ] = 1'd0;
    assign memhint[669 ] = 1'd0;
    assign memhint[670 ] = 1'd0;
    assign memhint[671 ] = 1'd0;
    assign memhint[672 ] = 1'd0;
    assign memhint[673 ] = 1'd0;
    assign memhint[674 ] = 1'd0;
    assign memhint[675 ] = 1'd1;
    assign memhint[676 ] = 1'd1;
    assign memhint[677 ] = 1'd1;
    assign memhint[678 ] = 1'd1;
    assign memhint[679 ] = 1'd1;
    assign memhint[680 ] = 1'd1;
    assign memhint[681 ] = 1'd1;
    assign memhint[682 ] = 1'd1;
    assign memhint[683 ] = 1'd1;
    assign memhint[684 ] = 1'd1;
    assign memhint[685 ] = 1'd1;
    assign memhint[686 ] = 1'd1;
    assign memhint[687 ] = 1'd0;
    assign memhint[688 ] = 1'd0;
    assign memhint[689 ] = 1'd0;
    assign memhint[690 ] = 1'd0;
    assign memhint[691 ] = 1'd0;
    assign memhint[692 ] = 1'd0;
    assign memhint[693 ] = 1'd0;
    assign memhint[694 ] = 1'd1;
    assign memhint[695 ] = 1'd1;
    assign memhint[696 ] = 1'd0;
    assign memhint[697 ] = 1'd0;
    assign memhint[698 ] = 1'd0;
    assign memhint[699 ] = 1'd0;
    assign memhint[700 ] = 1'd0;
    assign memhint[701 ] = 1'd0;
    assign memhint[702 ] = 1'd0;
    assign memhint[703 ] = 1'd0;
    assign memhint[704 ] = 1'd0;
    assign memhint[705 ] = 1'd0;
    assign memhint[706 ] = 1'd0;
    assign memhint[707 ] = 1'd0;
    assign memhint[708 ] = 1'd0;
    assign memhint[709 ] = 1'd0;
    assign memhint[710 ] = 1'd0;
    assign memhint[711 ] = 1'd0;
    assign memhint[712 ] = 1'd0;
    assign memhint[713 ] = 1'd0;
    assign memhint[714 ] = 1'd0;
    assign memhint[715 ] = 1'd0;
    assign memhint[716 ] = 1'd1;
    assign memhint[717 ] = 1'd1;
    assign memhint[718 ] = 1'd1;
    assign memhint[719 ] = 1'd0;
    assign memhint[720 ] = 1'd0;
    assign memhint[721 ] = 1'd0;
    assign memhint[722 ] = 1'd0;
    assign memhint[723 ] = 1'd0;
    assign memhint[724 ] = 1'd0;
    assign memhint[725 ] = 1'd0;
    assign memhint[726 ] = 1'd0;
    assign memhint[727 ] = 1'd0;
    assign memhint[728 ] = 1'd0;
    assign memhint[729 ] = 1'd0;
    assign memhint[730 ] = 1'd0;
    assign memhint[731 ] = 1'd1;
    assign memhint[732 ] = 1'd1;
    assign memhint[733 ] = 1'd0;
    assign memhint[734 ] = 1'd0;
    assign memhint[735 ] = 1'd0;
    assign memhint[736 ] = 1'd0;
    assign memhint[737 ] = 1'd0;
    assign memhint[738 ] = 1'd0;
    assign memhint[739 ] = 1'd0;
    assign memhint[740 ] = 1'd0;
    assign memhint[741 ] = 1'd0;
    assign memhint[742 ] = 1'd0;
    assign memhint[743 ] = 1'd1;
    assign memhint[744 ] = 1'd1;
    assign memhint[745 ] = 1'd0;
    assign memhint[746 ] = 1'd0;
    assign memhint[747 ] = 1'd0;
    assign memhint[748 ] = 1'd1;
    assign memhint[749 ] = 1'd1;
    assign memhint[750 ] = 1'd0;
    assign memhint[751 ] = 1'd0;
    assign memhint[752 ] = 1'd0;
    assign memhint[753 ] = 1'd0;
    assign memhint[754 ] = 1'd0;
    assign memhint[755 ] = 1'd1;
    assign memhint[756 ] = 1'd1;
    assign memhint[757 ] = 1'd1;
    assign memhint[758 ] = 1'd0;
    assign memhint[759 ] = 1'd0;
    assign memhint[760 ] = 1'd0;
    assign memhint[761 ] = 1'd0;
    assign memhint[762 ] = 1'd0;
    assign memhint[763 ] = 1'd0;
    assign memhint[764 ] = 1'd1;
    assign memhint[765 ] = 1'd1;
    assign memhint[766 ] = 1'd0;
    assign memhint[767 ] = 1'd0;
    assign memhint[768 ] = 1'd0;
    assign memhint[769 ] = 1'd0;
    assign memhint[770 ] = 1'd0;
    assign memhint[771 ] = 1'd0;
    assign memhint[772 ] = 1'd0;
    assign memhint[773 ] = 1'd0;
    assign memhint[774 ] = 1'd0;
    assign memhint[775 ] = 1'd0;
    assign memhint[776 ] = 1'd0;
    assign memhint[777 ] = 1'd0;
    assign memhint[778 ] = 1'd0;
    assign memhint[779 ] = 1'd0;
    assign memhint[780 ] = 1'd0;
    assign memhint[781 ] = 1'd1;
    assign memhint[782 ] = 1'd1;
    assign memhint[783 ] = 1'd0;
    assign memhint[784 ] = 1'd0;
    assign memhint[785 ] = 1'd0;
    assign memhint[786 ] = 1'd0;
    assign memhint[787 ] = 1'd0;
    assign memhint[788 ] = 1'd0;
    assign memhint[789 ] = 1'd0;
    assign memhint[790 ] = 1'd0;
    assign memhint[791 ] = 1'd0;
    assign memhint[792 ] = 1'd0;
    assign memhint[793 ] = 1'd0;
    assign memhint[794 ] = 1'd0;
    assign memhint[795 ] = 1'd0;
    assign memhint[796 ] = 1'd1;
    assign memhint[797 ] = 1'd1;
    assign memhint[798 ] = 1'd0;
    assign memhint[799 ] = 1'd0;
    assign memhint[800 ] = 1'd0;
    assign memhint[801 ] = 1'd0;
    assign memhint[802 ] = 1'd0;
    assign memhint[803 ] = 1'd0;
    assign memhint[804 ] = 1'd0;
    assign memhint[805 ] = 1'd0;
    assign memhint[806 ] = 1'd0;
    assign memhint[807 ] = 1'd0;
    assign memhint[808 ] = 1'd0;
    assign memhint[809 ] = 1'd0;
    assign memhint[810 ] = 1'd0;
    assign memhint[811 ] = 1'd0;
    assign memhint[812 ] = 1'd0;
    assign memhint[813 ] = 1'd0;
    assign memhint[814 ] = 1'd0;
    assign memhint[815 ] = 1'd0;
    assign memhint[816 ] = 1'd1;
    assign memhint[817 ] = 1'd1;
    assign memhint[818 ] = 1'd1;
    assign memhint[819 ] = 1'd1;
    assign memhint[820 ] = 1'd1;
    assign memhint[821 ] = 1'd0;
    assign memhint[822 ] = 1'd0;
    assign memhint[823 ] = 1'd0;
    assign memhint[824 ] = 1'd0;
    assign memhint[825 ] = 1'd0;
    assign memhint[826 ] = 1'd0;
    assign memhint[827 ] = 1'd1;
    assign memhint[828 ] = 1'd1;
    assign memhint[829 ] = 1'd1;
    assign memhint[830 ] = 1'd1;
    assign memhint[831 ] = 1'd1;
    assign memhint[832 ] = 1'd0;
    assign memhint[833 ] = 1'd0;
    assign memhint[834 ] = 1'd0;
    assign memhint[835 ] = 1'd0;
    assign memhint[836 ] = 1'd0;
    assign memhint[837 ] = 1'd0;
    assign memhint[838 ] = 1'd0;
    assign memhint[839 ] = 1'd0;
    assign memhint[840 ] = 1'd0;
    assign memhint[841 ] = 1'd1;
    assign memhint[842 ] = 1'd1;
    assign memhint[843 ] = 1'd0;
    assign memhint[844 ] = 1'd0;
    assign memhint[845 ] = 1'd0;
    assign memhint[846 ] = 1'd0;
    assign memhint[847 ] = 1'd0;
    assign memhint[848 ] = 1'd0;
    assign memhint[849 ] = 1'd0;
    assign memhint[850 ] = 1'd0;
    assign memhint[851 ] = 1'd0;
    assign memhint[852 ] = 1'd0;
    assign memhint[853 ] = 1'd0;
    assign memhint[854 ] = 1'd0;
    assign memhint[855 ] = 1'd0;
    assign memhint[856 ] = 1'd0;
    assign memhint[857 ] = 1'd0;
    assign memhint[858 ] = 1'd0;
    assign memhint[859 ] = 1'd0;
    assign memhint[860 ] = 1'd0;
    assign memhint[861 ] = 1'd0;
    assign memhint[862 ] = 1'd0;
    assign memhint[863 ] = 1'd0;
    assign memhint[864 ] = 1'd0;
    assign memhint[865 ] = 1'd0;
    assign memhint[866 ] = 1'd0;
    assign memhint[867 ] = 1'd0;
    assign memhint[868 ] = 1'd1;
    assign memhint[869 ] = 1'd1;
    assign memhint[870 ] = 1'd1;
    assign memhint[871 ] = 1'd0;
    assign memhint[872 ] = 1'd0;
    assign memhint[873 ] = 1'd0;
    assign memhint[874 ] = 1'd0;
    assign memhint[875 ] = 1'd0;
    assign memhint[876 ] = 1'd0;
    assign memhint[877 ] = 1'd0;
    assign memhint[878 ] = 1'd0;
    assign memhint[879 ] = 1'd0;
    assign memhint[880 ] = 1'd0;
    assign memhint[881 ] = 1'd0;
    assign memhint[882 ] = 1'd0;
    assign memhint[883 ] = 1'd0;
    assign memhint[884 ] = 1'd0;
    assign memhint[885 ] = 1'd0;
    assign memhint[886 ] = 1'd0;
    assign memhint[887 ] = 1'd0;
    assign memhint[888 ] = 1'd0;
    assign memhint[889 ] = 1'd0;
    assign memhint[890 ] = 1'd0;
    assign memhint[891 ] = 1'd0;
    assign memhint[892 ] = 1'd0;
    assign memhint[893 ] = 1'd1;
    assign memhint[894 ] = 1'd1;
    assign memhint[895 ] = 1'd0;
    assign memhint[896 ] = 1'd0;
    assign memhint[897 ] = 1'd0;
    assign memhint[898 ] = 1'd0;
    assign memhint[899 ] = 1'd0;
    assign memhint[900 ] = 1'd1;
    assign memhint[901 ] = 1'd1;
    assign memhint[902 ] = 1'd1;
    assign memhint[903 ] = 1'd0;
    assign memhint[904 ] = 1'd0;
    assign memhint[905 ] = 1'd0;
    assign memhint[906 ] = 1'd0;
    assign memhint[907 ] = 1'd0;
    assign memhint[908 ] = 1'd0;
    assign memhint[909 ] = 1'd0;
    assign memhint[910 ] = 1'd0;
    assign memhint[911 ] = 1'd0;
    assign memhint[912 ] = 1'd1;
    assign memhint[913 ] = 1'd1;
    assign memhint[914 ] = 1'd1;
    assign memhint[915 ] = 1'd1;
    assign memhint[916 ] = 1'd1;
    assign memhint[917 ] = 1'd0;
    assign memhint[918 ] = 1'd0;
    assign memhint[919 ] = 1'd0;
    assign memhint[920 ] = 1'd0;
    assign memhint[921 ] = 1'd0;
    assign memhint[922 ] = 1'd0;
    assign memhint[923 ] = 1'd1;
    assign memhint[924 ] = 1'd1;
    assign memhint[925 ] = 1'd1;
    assign memhint[926 ] = 1'd1;
    assign memhint[927 ] = 1'd1;
    assign memhint[928 ] = 1'd0;
    assign memhint[929 ] = 1'd0;
    assign memhint[930 ] = 1'd0;
    assign memhint[931 ] = 1'd0;
    assign memhint[932 ] = 1'd0;
    assign memhint[933 ] = 1'd0;
    assign memhint[934 ] = 1'd0;
    assign memhint[935 ] = 1'd0;
    assign memhint[936 ] = 1'd0;
    assign memhint[937 ] = 1'd1;
    assign memhint[938 ] = 1'd1;
    assign memhint[939 ] = 1'd1;
    assign memhint[940 ] = 1'd0;
    assign memhint[941 ] = 1'd0;
    assign memhint[942 ] = 1'd0;
    assign memhint[943 ] = 1'd0;
    assign memhint[944 ] = 1'd0;
    assign memhint[945 ] = 1'd0;
    assign memhint[946 ] = 1'd0;
    assign memhint[947 ] = 1'd0;
    assign memhint[948 ] = 1'd0;
    assign memhint[949 ] = 1'd0;
    assign memhint[950 ] = 1'd0;
    assign memhint[951 ] = 1'd0;
    assign memhint[952 ] = 1'd0;
    assign memhint[953 ] = 1'd1;
    assign memhint[954 ] = 1'd1;
    assign memhint[955 ] = 1'd0;
    assign memhint[956 ] = 1'd0;
    assign memhint[957 ] = 1'd0;
    assign memhint[958 ] = 1'd0;
    assign memhint[959 ] = 1'd0;
    assign memhint[960 ] = 1'd0;
    assign memhint[961 ] = 1'd0;
    assign memhint[962 ] = 1'd0;
    assign memhint[963 ] = 1'd0;
    assign memhint[964 ] = 1'd0;
    assign memhint[965 ] = 1'd1;
    assign memhint[966 ] = 1'd1;
    assign memhint[967 ] = 1'd1;
    assign memhint[968 ] = 1'd1;
    assign memhint[969 ] = 1'd0;
    assign memhint[970 ] = 1'd0;
    assign memhint[971 ] = 1'd0;
    assign memhint[972 ] = 1'd0;
    assign memhint[973 ] = 1'd0;
    assign memhint[974 ] = 1'd0;
    assign memhint[975 ] = 1'd0;
    assign memhint[976 ] = 1'd1;
    assign memhint[977 ] = 1'd1;
    assign memhint[978 ] = 1'd1;
    assign memhint[979 ] = 1'd1;
    assign memhint[980 ] = 1'd1;
    assign memhint[981 ] = 1'd0;
    assign memhint[982 ] = 1'd0;
    assign memhint[983 ] = 1'd0;
    assign memhint[984 ] = 1'd0;
    assign memhint[985 ] = 1'd0;
    assign memhint[986 ] = 1'd0;
    assign memhint[987 ] = 1'd0;
    assign memhint[988 ] = 1'd0;
    assign memhint[989 ] = 1'd0;
    assign memhint[990 ] = 1'd0;
    assign memhint[991 ] = 1'd0;
    assign memhint[992 ] = 1'd0;
    assign memhint[993 ] = 1'd0;
    assign memhint[994 ] = 1'd0;
    assign memhint[995 ] = 1'd0;
    assign memhint[996 ] = 1'd0;
    assign memhint[997 ] = 1'd0;
    assign memhint[998 ] = 1'd0;
    assign memhint[999 ] = 1'd0;
    assign memhint[1000] = 1'd1;
    assign memhint[1001] = 1'd1;
    assign memhint[1002] = 1'd0;
    assign memhint[1003] = 1'd0;
    assign memhint[1004] = 1'd0;
    assign memhint[1005] = 1'd0;
    assign memhint[1006] = 1'd0;
    assign memhint[1007] = 1'd0;
    assign memhint[1008] = 1'd0;
    assign memhint[1009] = 1'd0;
    assign memhint[1010] = 1'd0;
    assign memhint[1011] = 1'd0;
    assign memhint[1012] = 1'd0;
    assign memhint[1013] = 1'd0;
    assign memhint[1014] = 1'd1;
    assign memhint[1015] = 1'd1;
    assign memhint[1016] = 1'd1;
    assign memhint[1017] = 1'd1;
    assign memhint[1018] = 1'd1;
    assign memhint[1019] = 1'd0;
    assign memhint[1020] = 1'd0;
    assign memhint[1021] = 1'd0;
    assign memhint[1022] = 1'd0;
    assign memhint[1023] = 1'd0;
    assign memhint[1024] = 1'd0;
    assign memhint[1025] = 1'd1;
    assign memhint[1026] = 1'd1;
    assign memhint[1027] = 1'd1;
    assign memhint[1028] = 1'd1;
    assign memhint[1029] = 1'd1;
    assign memhint[1030] = 1'd0;
    assign memhint[1031] = 1'd0;
    assign memhint[1032] = 1'd0;
    assign memhint[1033] = 1'd0;
    assign memhint[1034] = 1'd0;
    assign memhint[1035] = 1'd0;
    assign memhint[1036] = 1'd0;
    assign memhint[1037] = 1'd0;
    assign memhint[1038] = 1'd0;
    assign memhint[1039] = 1'd0;
    assign memhint[1040] = 1'd0;
    assign memhint[1041] = 1'd0;
    assign memhint[1042] = 1'd0;
    assign memhint[1043] = 1'd0;
    assign memhint[1044] = 1'd0;
    assign memhint[1045] = 1'd0;
    assign memhint[1046] = 1'd0;
    assign memhint[1047] = 1'd0;
    assign memhint[1048] = 1'd1;
    assign memhint[1049] = 1'd1;
    assign memhint[1050] = 1'd0;
    assign memhint[1051] = 1'd0;
    assign memhint[1052] = 1'd0;
    assign memhint[1053] = 1'd0;
    assign memhint[1054] = 1'd0;
    assign memhint[1055] = 1'd0;
    assign memhint[1056] = 1'd0;
    assign memhint[1057] = 1'd0;
    assign memhint[1058] = 1'd1;
    assign memhint[1059] = 1'd1;
    assign memhint[1060] = 1'd1;
    assign memhint[1061] = 1'd0;
    assign memhint[1062] = 1'd0;
    assign memhint[1063] = 1'd0;
    assign memhint[1064] = 1'd0;
    assign memhint[1065] = 1'd0;
    assign memhint[1066] = 1'd0;
    assign memhint[1067] = 1'd1;
    assign memhint[1068] = 1'd1;
    assign memhint[1069] = 1'd0;
    assign memhint[1070] = 1'd0;
    assign memhint[1071] = 1'd0;
    assign memhint[1072] = 1'd0;
    assign memhint[1073] = 1'd0;
    assign memhint[1074] = 1'd0;
    assign memhint[1075] = 1'd0;
    assign memhint[1076] = 1'd0;
    assign memhint[1077] = 1'd0;
    assign memhint[1078] = 1'd0;
    assign memhint[1079] = 1'd0;
    assign memhint[1080] = 1'd0;
    assign memhint[1081] = 1'd0;
    assign memhint[1082] = 1'd0;
    assign memhint[1083] = 1'd0;
    assign memhint[1084] = 1'd0;
    assign memhint[1085] = 1'd0;
    assign memhint[1086] = 1'd0;
    assign memhint[1087] = 1'd0;
    assign memhint[1088] = 1'd0;
    assign memhint[1089] = 1'd1;
    assign memhint[1090] = 1'd1;
    assign memhint[1091] = 1'd1;
    assign memhint[1092] = 1'd0;
    assign memhint[1093] = 1'd0;
    assign memhint[1094] = 1'd0;
    assign memhint[1095] = 1'd0;
    assign memhint[1096] = 1'd0;
    assign memhint[1097] = 1'd0;
    assign memhint[1098] = 1'd0;
    assign memhint[1099] = 1'd0;
    assign memhint[1100] = 1'd0;
    assign memhint[1101] = 1'd0;
    assign memhint[1102] = 1'd0;
    assign memhint[1103] = 1'd0;
    assign memhint[1104] = 1'd1;
    assign memhint[1105] = 1'd1;
    assign memhint[1106] = 1'd1;
    assign memhint[1107] = 1'd0;
    assign memhint[1108] = 1'd0;
    assign memhint[1109] = 1'd0;
    assign memhint[1110] = 1'd0;
    assign memhint[1111] = 1'd0;
    assign memhint[1112] = 1'd0;
    assign memhint[1113] = 1'd0;
    assign memhint[1114] = 1'd0;
    assign memhint[1115] = 1'd1;
    assign memhint[1116] = 1'd1;
    assign memhint[1117] = 1'd1;
    assign memhint[1118] = 1'd0;
    assign memhint[1119] = 1'd0;
    assign memhint[1120] = 1'd1;
    assign memhint[1121] = 1'd1;
    assign memhint[1122] = 1'd0;
    assign memhint[1123] = 1'd0;
    assign memhint[1124] = 1'd0;
    assign memhint[1125] = 1'd0;
    assign memhint[1126] = 1'd0;
    assign memhint[1127] = 1'd0;
    assign memhint[1128] = 1'd0;
    assign memhint[1129] = 1'd1;
    assign memhint[1130] = 1'd1;
    assign memhint[1131] = 1'd1;
    assign memhint[1132] = 1'd0;
    assign memhint[1133] = 1'd0;
    assign memhint[1134] = 1'd0;
    assign memhint[1135] = 1'd0;
    assign memhint[1136] = 1'd0;
    assign memhint[1137] = 1'd1;
    assign memhint[1138] = 1'd1;
    assign memhint[1139] = 1'd0;
    assign memhint[1140] = 1'd0;
    assign memhint[1141] = 1'd0;
    assign memhint[1142] = 1'd0;
    assign memhint[1143] = 1'd0;
    assign memhint[1144] = 1'd0;
    assign memhint[1145] = 1'd0;
    assign memhint[1146] = 1'd0;
    assign memhint[1147] = 1'd0;
    assign memhint[1148] = 1'd0;
    assign memhint[1149] = 1'd0;
    assign memhint[1150] = 1'd0;
    assign memhint[1151] = 1'd0;
    assign memhint[1152] = 1'd0;
    assign memhint[1153] = 1'd0;
    assign memhint[1154] = 1'd1;
    assign memhint[1155] = 1'd1;
    assign memhint[1156] = 1'd0;
    assign memhint[1157] = 1'd0;
    assign memhint[1158] = 1'd0;
    assign memhint[1159] = 1'd0;
    assign memhint[1160] = 1'd0;
    assign memhint[1161] = 1'd0;
    assign memhint[1162] = 1'd0;
    assign memhint[1163] = 1'd0;
    assign memhint[1164] = 1'd0;
    assign memhint[1165] = 1'd0;
    assign memhint[1166] = 1'd0;
    assign memhint[1167] = 1'd0;
    assign memhint[1168] = 1'd0;
    assign memhint[1169] = 1'd1;
    assign memhint[1170] = 1'd1;
    assign memhint[1171] = 1'd0;
    assign memhint[1172] = 1'd0;
    assign memhint[1173] = 1'd0;
    assign memhint[1174] = 1'd0;
    assign memhint[1175] = 1'd0;
    assign memhint[1176] = 1'd0;
    assign memhint[1177] = 1'd0;
    assign memhint[1178] = 1'd0;
    assign memhint[1179] = 1'd0;
    assign memhint[1180] = 1'd0;
    assign memhint[1181] = 1'd0;
    assign memhint[1182] = 1'd0;
    assign memhint[1183] = 1'd0;
    assign memhint[1184] = 1'd0;
    assign memhint[1185] = 1'd0;
    assign memhint[1186] = 1'd0;
    assign memhint[1187] = 1'd0;
    assign memhint[1188] = 1'd1;
    assign memhint[1189] = 1'd1;
    assign memhint[1190] = 1'd1;
    assign memhint[1191] = 1'd1;
    assign memhint[1192] = 1'd0;
    assign memhint[1193] = 1'd0;
    assign memhint[1194] = 1'd0;
    assign memhint[1195] = 1'd0;
    assign memhint[1196] = 1'd0;
    assign memhint[1197] = 1'd0;
    assign memhint[1198] = 1'd0;
    assign memhint[1199] = 1'd0;
    assign memhint[1200] = 1'd0;
    assign memhint[1201] = 1'd0;
    assign memhint[1202] = 1'd1;
    assign memhint[1203] = 1'd1;
    assign memhint[1204] = 1'd1;
    assign memhint[1205] = 1'd1;
    assign memhint[1206] = 1'd0;
    assign memhint[1207] = 1'd0;
    assign memhint[1208] = 1'd0;
    assign memhint[1209] = 1'd0;
    assign memhint[1210] = 1'd0;
    assign memhint[1211] = 1'd0;
    assign memhint[1212] = 1'd0;
    assign memhint[1213] = 1'd0;
    assign memhint[1214] = 1'd1;
    assign memhint[1215] = 1'd1;
    assign memhint[1216] = 1'd0;
    assign memhint[1217] = 1'd0;
    assign memhint[1218] = 1'd0;
    assign memhint[1219] = 1'd0;
    assign memhint[1220] = 1'd0;
    assign memhint[1221] = 1'd0;
    assign memhint[1222] = 1'd0;
    assign memhint[1223] = 1'd0;
    assign memhint[1224] = 1'd0;
    assign memhint[1225] = 1'd0;
    assign memhint[1226] = 1'd0;
    assign memhint[1227] = 1'd0;
    assign memhint[1228] = 1'd0;
    assign memhint[1229] = 1'd0;
    assign memhint[1230] = 1'd0;
    assign memhint[1231] = 1'd0;
    assign memhint[1232] = 1'd0;
    assign memhint[1233] = 1'd0;
    assign memhint[1234] = 1'd0;
    assign memhint[1235] = 1'd0;
    assign memhint[1236] = 1'd0;
    assign memhint[1237] = 1'd0;
    assign memhint[1238] = 1'd0;
    assign memhint[1239] = 1'd0;
    assign memhint[1240] = 1'd1;
    assign memhint[1241] = 1'd1;
    assign memhint[1242] = 1'd1;
    assign memhint[1243] = 1'd1;
    assign memhint[1244] = 1'd1;
    assign memhint[1245] = 1'd0;
    assign memhint[1246] = 1'd0;
    assign memhint[1247] = 1'd0;
    assign memhint[1248] = 1'd0;
    assign memhint[1249] = 1'd0;
    assign memhint[1250] = 1'd0;
    assign memhint[1251] = 1'd0;
    assign memhint[1252] = 1'd0;
    assign memhint[1253] = 1'd0;
    assign memhint[1254] = 1'd0;
    assign memhint[1255] = 1'd0;
    assign memhint[1256] = 1'd0;
    assign memhint[1257] = 1'd0;
    assign memhint[1258] = 1'd0;
    assign memhint[1259] = 1'd0;
    assign memhint[1260] = 1'd0;
    assign memhint[1261] = 1'd0;
    assign memhint[1262] = 1'd0;
    assign memhint[1263] = 1'd0;
    assign memhint[1264] = 1'd0;
    assign memhint[1265] = 1'd1;
    assign memhint[1266] = 1'd1;
    assign memhint[1267] = 1'd0;
    assign memhint[1268] = 1'd0;
    assign memhint[1269] = 1'd0;
    assign memhint[1270] = 1'd0;
    assign memhint[1271] = 1'd0;
    assign memhint[1272] = 1'd0;
    assign memhint[1273] = 1'd0;
    assign memhint[1274] = 1'd1;
    assign memhint[1275] = 1'd1;
    assign memhint[1276] = 1'd1;
    assign memhint[1277] = 1'd0;
    assign memhint[1278] = 1'd0;
    assign memhint[1279] = 1'd0;
    assign memhint[1280] = 1'd0;
    assign memhint[1281] = 1'd0;
    assign memhint[1282] = 1'd0;
    assign memhint[1283] = 1'd0;
    assign memhint[1284] = 1'd1;
    assign memhint[1285] = 1'd1;
    assign memhint[1286] = 1'd1;
    assign memhint[1287] = 1'd1;
    assign memhint[1288] = 1'd0;
    assign memhint[1289] = 1'd0;
    assign memhint[1290] = 1'd0;
    assign memhint[1291] = 1'd0;
    assign memhint[1292] = 1'd0;
    assign memhint[1293] = 1'd0;
    assign memhint[1294] = 1'd0;
    assign memhint[1295] = 1'd0;
    assign memhint[1296] = 1'd0;
    assign memhint[1297] = 1'd0;
    assign memhint[1298] = 1'd1;
    assign memhint[1299] = 1'd1;
    assign memhint[1300] = 1'd1;
    assign memhint[1301] = 1'd1;
    assign memhint[1302] = 1'd0;
    assign memhint[1303] = 1'd0;
    assign memhint[1304] = 1'd0;
    assign memhint[1305] = 1'd0;
    assign memhint[1306] = 1'd0;
    assign memhint[1307] = 1'd0;
    assign memhint[1308] = 1'd0;
    assign memhint[1309] = 1'd0;
    assign memhint[1310] = 1'd1;
    assign memhint[1311] = 1'd1;
    assign memhint[1312] = 1'd1;
    assign memhint[1313] = 1'd0;
    assign memhint[1314] = 1'd0;
    assign memhint[1315] = 1'd0;
    assign memhint[1316] = 1'd0;
    assign memhint[1317] = 1'd0;
    assign memhint[1318] = 1'd0;
    assign memhint[1319] = 1'd0;
    assign memhint[1320] = 1'd0;
    assign memhint[1321] = 1'd0;
    assign memhint[1322] = 1'd0;
    assign memhint[1323] = 1'd0;
    assign memhint[1324] = 1'd0;
    assign memhint[1325] = 1'd0;
    assign memhint[1326] = 1'd1;
    assign memhint[1327] = 1'd1;
    assign memhint[1328] = 1'd0;
    assign memhint[1329] = 1'd0;
    assign memhint[1330] = 1'd0;
    assign memhint[1331] = 1'd0;
    assign memhint[1332] = 1'd0;
    assign memhint[1333] = 1'd0;
    assign memhint[1334] = 1'd0;
    assign memhint[1335] = 1'd0;
    assign memhint[1336] = 1'd1;
    assign memhint[1337] = 1'd1;
    assign memhint[1338] = 1'd1;
    assign memhint[1339] = 1'd1;
    assign memhint[1340] = 1'd0;
    assign memhint[1341] = 1'd0;
    assign memhint[1342] = 1'd0;
    assign memhint[1343] = 1'd0;
    assign memhint[1344] = 1'd0;
    assign memhint[1345] = 1'd0;
    assign memhint[1346] = 1'd0;
    assign memhint[1347] = 1'd0;
    assign memhint[1348] = 1'd0;
    assign memhint[1349] = 1'd0;
    assign memhint[1350] = 1'd0;
    assign memhint[1351] = 1'd1;
    assign memhint[1352] = 1'd1;
    assign memhint[1353] = 1'd1;
    assign memhint[1354] = 1'd1;
    assign memhint[1355] = 1'd0;
    assign memhint[1356] = 1'd0;
    assign memhint[1357] = 1'd0;
    assign memhint[1358] = 1'd0;
    assign memhint[1359] = 1'd0;
    assign memhint[1360] = 1'd0;
    assign memhint[1361] = 1'd0;
    assign memhint[1362] = 1'd0;
    assign memhint[1363] = 1'd0;
    assign memhint[1364] = 1'd0;
    assign memhint[1365] = 1'd0;
    assign memhint[1366] = 1'd0;
    assign memhint[1367] = 1'd0;
    assign memhint[1368] = 1'd0;
    assign memhint[1369] = 1'd0;
    assign memhint[1370] = 1'd0;
    assign memhint[1371] = 1'd0;
    assign memhint[1372] = 1'd0;
    assign memhint[1373] = 1'd1;
    assign memhint[1374] = 1'd1;
    assign memhint[1375] = 1'd0;
    assign memhint[1376] = 1'd0;
    assign memhint[1377] = 1'd0;
    assign memhint[1378] = 1'd0;
    assign memhint[1379] = 1'd0;
    assign memhint[1380] = 1'd0;
    assign memhint[1381] = 1'd0;
    assign memhint[1382] = 1'd0;
    assign memhint[1383] = 1'd0;
    assign memhint[1384] = 1'd0;
    assign memhint[1385] = 1'd0;
    assign memhint[1386] = 1'd1;
    assign memhint[1387] = 1'd1;
    assign memhint[1388] = 1'd1;
    assign memhint[1389] = 1'd1;
    assign memhint[1390] = 1'd0;
    assign memhint[1391] = 1'd0;
    assign memhint[1392] = 1'd0;
    assign memhint[1393] = 1'd0;
    assign memhint[1394] = 1'd0;
    assign memhint[1395] = 1'd0;
    assign memhint[1396] = 1'd0;
    assign memhint[1397] = 1'd0;
    assign memhint[1398] = 1'd0;
    assign memhint[1399] = 1'd0;
    assign memhint[1400] = 1'd1;
    assign memhint[1401] = 1'd1;
    assign memhint[1402] = 1'd1;
    assign memhint[1403] = 1'd1;
    assign memhint[1404] = 1'd0;
    assign memhint[1405] = 1'd0;
    assign memhint[1406] = 1'd0;
    assign memhint[1407] = 1'd0;
    assign memhint[1408] = 1'd0;
    assign memhint[1409] = 1'd0;
    assign memhint[1410] = 1'd0;
    assign memhint[1411] = 1'd0;
    assign memhint[1412] = 1'd0;
    assign memhint[1413] = 1'd0;
    assign memhint[1414] = 1'd0;
    assign memhint[1415] = 1'd0;
    assign memhint[1416] = 1'd0;
    assign memhint[1417] = 1'd0;
    assign memhint[1418] = 1'd0;
    assign memhint[1419] = 1'd0;
    assign memhint[1420] = 1'd0;
    assign memhint[1421] = 1'd1;
    assign memhint[1422] = 1'd1;
    assign memhint[1423] = 1'd0;
    assign memhint[1424] = 1'd0;
    assign memhint[1425] = 1'd0;
    assign memhint[1426] = 1'd0;
    assign memhint[1427] = 1'd0;
    assign memhint[1428] = 1'd0;
    assign memhint[1429] = 1'd0;
    assign memhint[1430] = 1'd0;
    assign memhint[1431] = 1'd0;
    assign memhint[1432] = 1'd1;
    assign memhint[1433] = 1'd1;
    assign memhint[1434] = 1'd1;
    assign memhint[1435] = 1'd0;
    assign memhint[1436] = 1'd0;
    assign memhint[1437] = 1'd0;
    assign memhint[1438] = 1'd0;
    assign memhint[1439] = 1'd0;
    assign memhint[1440] = 1'd1;
    assign memhint[1441] = 1'd1;
    assign memhint[1442] = 1'd0;
    assign memhint[1443] = 1'd0;
    assign memhint[1444] = 1'd0;
    assign memhint[1445] = 1'd0;
    assign memhint[1446] = 1'd0;
    assign memhint[1447] = 1'd0;
    assign memhint[1448] = 1'd0;
    assign memhint[1449] = 1'd0;
    assign memhint[1450] = 1'd0;
    assign memhint[1451] = 1'd0;
    assign memhint[1452] = 1'd0;
    assign memhint[1453] = 1'd0;
    assign memhint[1454] = 1'd0;
    assign memhint[1455] = 1'd0;
    assign memhint[1456] = 1'd0;
    assign memhint[1457] = 1'd0;
    assign memhint[1458] = 1'd0;
    assign memhint[1459] = 1'd0;
    assign memhint[1460] = 1'd0;
    assign memhint[1461] = 1'd1;
    assign memhint[1462] = 1'd1;
    assign memhint[1463] = 1'd1;
    assign memhint[1464] = 1'd1;
    assign memhint[1465] = 1'd1;
    assign memhint[1466] = 1'd0;
    assign memhint[1467] = 1'd0;
    assign memhint[1468] = 1'd0;
    assign memhint[1469] = 1'd0;
    assign memhint[1470] = 1'd0;
    assign memhint[1471] = 1'd0;
    assign memhint[1472] = 1'd0;
    assign memhint[1473] = 1'd0;
    assign memhint[1474] = 1'd0;
    assign memhint[1475] = 1'd0;
    assign memhint[1476] = 1'd0;
    assign memhint[1477] = 1'd0;
    assign memhint[1478] = 1'd1;
    assign memhint[1479] = 1'd1;
    assign memhint[1480] = 1'd0;
    assign memhint[1481] = 1'd0;
    assign memhint[1482] = 1'd0;
    assign memhint[1483] = 1'd0;
    assign memhint[1484] = 1'd0;
    assign memhint[1485] = 1'd0;
    assign memhint[1486] = 1'd0;
    assign memhint[1487] = 1'd0;
    assign memhint[1488] = 1'd1;
    assign memhint[1489] = 1'd1;
    assign memhint[1490] = 1'd0;
    assign memhint[1491] = 1'd0;
    assign memhint[1492] = 1'd0;
    assign memhint[1493] = 1'd1;
    assign memhint[1494] = 1'd1;
    assign memhint[1495] = 1'd0;
    assign memhint[1496] = 1'd0;
    assign memhint[1497] = 1'd0;
    assign memhint[1498] = 1'd0;
    assign memhint[1499] = 1'd0;
    assign memhint[1500] = 1'd0;
    assign memhint[1501] = 1'd0;
    assign memhint[1502] = 1'd0;
    assign memhint[1503] = 1'd1;
    assign memhint[1504] = 1'd0;
    assign memhint[1505] = 1'd0;
    assign memhint[1506] = 1'd0;
    assign memhint[1507] = 1'd0;
    assign memhint[1508] = 1'd0;
    assign memhint[1509] = 1'd0;
    assign memhint[1510] = 1'd1;
    assign memhint[1511] = 1'd1;
    assign memhint[1512] = 1'd0;
    assign memhint[1513] = 1'd0;
    assign memhint[1514] = 1'd0;
    assign memhint[1515] = 1'd0;
    assign memhint[1516] = 1'd0;
    assign memhint[1517] = 1'd0;
    assign memhint[1518] = 1'd0;
    assign memhint[1519] = 1'd0;
    assign memhint[1520] = 1'd0;
    assign memhint[1521] = 1'd0;
    assign memhint[1522] = 1'd0;
    assign memhint[1523] = 1'd0;
    assign memhint[1524] = 1'd0;
    assign memhint[1525] = 1'd0;
    assign memhint[1526] = 1'd0;
    assign memhint[1527] = 1'd1;
    assign memhint[1528] = 1'd1;
    assign memhint[1529] = 1'd0;
    assign memhint[1530] = 1'd0;
    assign memhint[1531] = 1'd0;
    assign memhint[1532] = 1'd0;
    assign memhint[1533] = 1'd0;
    assign memhint[1534] = 1'd0;
    assign memhint[1535] = 1'd0;
    assign memhint[1536] = 1'd0;
    assign memhint[1537] = 1'd0;
    assign memhint[1538] = 1'd0;
    assign memhint[1539] = 1'd0;
    assign memhint[1540] = 1'd0;
    assign memhint[1541] = 1'd0;
    assign memhint[1542] = 1'd1;
    assign memhint[1543] = 1'd1;
    assign memhint[1544] = 1'd0;
    assign memhint[1545] = 1'd0;
    assign memhint[1546] = 1'd0;
    assign memhint[1547] = 1'd0;
    assign memhint[1548] = 1'd0;
    assign memhint[1549] = 1'd0;
    assign memhint[1550] = 1'd0;
    assign memhint[1551] = 1'd0;
    assign memhint[1552] = 1'd0;
    assign memhint[1553] = 1'd0;
    assign memhint[1554] = 1'd0;
    assign memhint[1555] = 1'd0;
    assign memhint[1556] = 1'd0;
    assign memhint[1557] = 1'd0;
    assign memhint[1558] = 1'd0;
    assign memhint[1559] = 1'd0;
    assign memhint[1560] = 1'd1;
    assign memhint[1561] = 1'd1;
    assign memhint[1562] = 1'd1;
    assign memhint[1563] = 1'd0;
    assign memhint[1564] = 1'd0;
    assign memhint[1565] = 1'd0;
    assign memhint[1566] = 1'd0;
    assign memhint[1567] = 1'd0;
    assign memhint[1568] = 1'd0;
    assign memhint[1569] = 1'd0;
    assign memhint[1570] = 1'd0;
    assign memhint[1571] = 1'd0;
    assign memhint[1572] = 1'd0;
    assign memhint[1573] = 1'd0;
    assign memhint[1574] = 1'd0;
    assign memhint[1575] = 1'd0;
    assign memhint[1576] = 1'd0;
    assign memhint[1577] = 1'd1;
    assign memhint[1578] = 1'd1;
    assign memhint[1579] = 1'd1;
    assign memhint[1580] = 1'd0;
    assign memhint[1581] = 1'd0;
    assign memhint[1582] = 1'd0;
    assign memhint[1583] = 1'd0;
    assign memhint[1584] = 1'd0;
    assign memhint[1585] = 1'd0;
    assign memhint[1586] = 1'd0;
    assign memhint[1587] = 1'd1;
    assign memhint[1588] = 1'd1;
    assign memhint[1589] = 1'd0;
    assign memhint[1590] = 1'd0;
    assign memhint[1591] = 1'd0;
    assign memhint[1592] = 1'd0;
    assign memhint[1593] = 1'd0;
    assign memhint[1594] = 1'd0;
    assign memhint[1595] = 1'd0;
    assign memhint[1596] = 1'd0;
    assign memhint[1597] = 1'd0;
    assign memhint[1598] = 1'd0;
    assign memhint[1599] = 1'd0;
    assign memhint[1600] = 1'd0;
    assign memhint[1601] = 1'd0;
    assign memhint[1602] = 1'd0;
    assign memhint[1603] = 1'd0;
    assign memhint[1604] = 1'd0;
    assign memhint[1605] = 1'd0;
    assign memhint[1606] = 1'd0;
    assign memhint[1607] = 1'd0;
    assign memhint[1608] = 1'd0;
    assign memhint[1609] = 1'd0;
    assign memhint[1610] = 1'd0;
    assign memhint[1611] = 1'd0;
    assign memhint[1612] = 1'd0;
    assign memhint[1613] = 1'd1;
    assign memhint[1614] = 1'd1;
    assign memhint[1615] = 1'd0;
    assign memhint[1616] = 1'd1;
    assign memhint[1617] = 1'd1;
    assign memhint[1618] = 1'd0;
    assign memhint[1619] = 1'd0;
    assign memhint[1620] = 1'd0;
    assign memhint[1621] = 1'd0;
    assign memhint[1622] = 1'd0;
    assign memhint[1623] = 1'd0;
    assign memhint[1624] = 1'd0;
    assign memhint[1625] = 1'd0;
    assign memhint[1626] = 1'd0;
    assign memhint[1627] = 1'd0;
    assign memhint[1628] = 1'd0;
    assign memhint[1629] = 1'd0;
    assign memhint[1630] = 1'd0;
    assign memhint[1631] = 1'd0;
    assign memhint[1632] = 1'd0;
    assign memhint[1633] = 1'd0;
    assign memhint[1634] = 1'd0;
    assign memhint[1635] = 1'd0;
    assign memhint[1636] = 1'd0;
    assign memhint[1637] = 1'd0;
    assign memhint[1638] = 1'd1;
    assign memhint[1639] = 1'd1;
    assign memhint[1640] = 1'd0;
    assign memhint[1641] = 1'd0;
    assign memhint[1642] = 1'd0;
    assign memhint[1643] = 1'd0;
    assign memhint[1644] = 1'd0;
    assign memhint[1645] = 1'd0;
    assign memhint[1646] = 1'd0;
    assign memhint[1647] = 1'd0;
    assign memhint[1648] = 1'd1;
    assign memhint[1649] = 1'd0;
    assign memhint[1650] = 1'd0;
    assign memhint[1651] = 1'd0;
    assign memhint[1652] = 1'd0;
    assign memhint[1653] = 1'd0;
    assign memhint[1654] = 1'd0;
    assign memhint[1655] = 1'd0;
    assign memhint[1656] = 1'd1;
    assign memhint[1657] = 1'd1;
    assign memhint[1658] = 1'd1;
    assign memhint[1659] = 1'd0;
    assign memhint[1660] = 1'd0;
    assign memhint[1661] = 1'd0;
    assign memhint[1662] = 1'd0;
    assign memhint[1663] = 1'd0;
    assign memhint[1664] = 1'd0;
    assign memhint[1665] = 1'd0;
    assign memhint[1666] = 1'd0;
    assign memhint[1667] = 1'd0;
    assign memhint[1668] = 1'd0;
    assign memhint[1669] = 1'd0;
    assign memhint[1670] = 1'd0;
    assign memhint[1671] = 1'd0;
    assign memhint[1672] = 1'd0;
    assign memhint[1673] = 1'd1;
    assign memhint[1674] = 1'd1;
    assign memhint[1675] = 1'd1;
    assign memhint[1676] = 1'd0;
    assign memhint[1677] = 1'd0;
    assign memhint[1678] = 1'd0;
    assign memhint[1679] = 1'd0;
    assign memhint[1680] = 1'd0;
    assign memhint[1681] = 1'd0;
    assign memhint[1682] = 1'd0;
    assign memhint[1683] = 1'd1;
    assign memhint[1684] = 1'd1;
    assign memhint[1685] = 1'd1;
    assign memhint[1686] = 1'd1;
    assign memhint[1687] = 1'd0;
    assign memhint[1688] = 1'd0;
    assign memhint[1689] = 1'd0;
    assign memhint[1690] = 1'd0;
    assign memhint[1691] = 1'd0;
    assign memhint[1692] = 1'd0;
    assign memhint[1693] = 1'd0;
    assign memhint[1694] = 1'd0;
    assign memhint[1695] = 1'd0;
    assign memhint[1696] = 1'd0;
    assign memhint[1697] = 1'd0;
    assign memhint[1698] = 1'd0;
    assign memhint[1699] = 1'd1;
    assign memhint[1700] = 1'd1;
    assign memhint[1701] = 1'd0;
    assign memhint[1702] = 1'd0;
    assign memhint[1703] = 1'd0;
    assign memhint[1704] = 1'd0;
    assign memhint[1705] = 1'd0;
    assign memhint[1706] = 1'd0;
    assign memhint[1707] = 1'd0;
    assign memhint[1708] = 1'd1;
    assign memhint[1709] = 1'd1;
    assign memhint[1710] = 1'd1;
    assign memhint[1711] = 1'd0;
    assign memhint[1712] = 1'd0;
    assign memhint[1713] = 1'd0;
    assign memhint[1714] = 1'd0;
    assign memhint[1715] = 1'd0;
    assign memhint[1716] = 1'd0;
    assign memhint[1717] = 1'd0;
    assign memhint[1718] = 1'd0;
    assign memhint[1719] = 1'd0;
    assign memhint[1720] = 1'd0;
    assign memhint[1721] = 1'd0;
    assign memhint[1722] = 1'd0;
    assign memhint[1723] = 1'd0;
    assign memhint[1724] = 1'd0;
    assign memhint[1725] = 1'd1;
    assign memhint[1726] = 1'd1;
    assign memhint[1727] = 1'd1;
    assign memhint[1728] = 1'd1;
    assign memhint[1729] = 1'd0;
    assign memhint[1730] = 1'd0;
    assign memhint[1731] = 1'd0;
    assign memhint[1732] = 1'd0;
    assign memhint[1733] = 1'd0;
    assign memhint[1734] = 1'd0;
    assign memhint[1735] = 1'd0;
    assign memhint[1736] = 1'd0;
    assign memhint[1737] = 1'd0;
    assign memhint[1738] = 1'd0;
    assign memhint[1739] = 1'd0;
    assign memhint[1740] = 1'd0;
    assign memhint[1741] = 1'd0;
    assign memhint[1742] = 1'd0;
    assign memhint[1743] = 1'd0;
    assign memhint[1744] = 1'd0;
    assign memhint[1745] = 1'd0;
    assign memhint[1746] = 1'd1;
    assign memhint[1747] = 1'd1;
    assign memhint[1748] = 1'd0;
    assign memhint[1749] = 1'd0;
    assign memhint[1750] = 1'd0;
    assign memhint[1751] = 1'd0;
    assign memhint[1752] = 1'd0;
    assign memhint[1753] = 1'd0;
    assign memhint[1754] = 1'd0;
    assign memhint[1755] = 1'd0;
    assign memhint[1756] = 1'd0;
    assign memhint[1757] = 1'd0;
    assign memhint[1758] = 1'd1;
    assign memhint[1759] = 1'd1;
    assign memhint[1760] = 1'd1;
    assign memhint[1761] = 1'd0;
    assign memhint[1762] = 1'd0;
    assign memhint[1763] = 1'd0;
    assign memhint[1764] = 1'd0;
    assign memhint[1765] = 1'd0;
    assign memhint[1766] = 1'd0;
    assign memhint[1767] = 1'd0;
    assign memhint[1768] = 1'd0;
    assign memhint[1769] = 1'd0;
    assign memhint[1770] = 1'd0;
    assign memhint[1771] = 1'd0;
    assign memhint[1772] = 1'd0;
    assign memhint[1773] = 1'd0;
    assign memhint[1774] = 1'd0;
    assign memhint[1775] = 1'd1;
    assign memhint[1776] = 1'd1;
    assign memhint[1777] = 1'd1;
    assign memhint[1778] = 1'd0;
    assign memhint[1779] = 1'd0;
    assign memhint[1780] = 1'd0;
    assign memhint[1781] = 1'd0;
    assign memhint[1782] = 1'd0;
    assign memhint[1783] = 1'd0;
    assign memhint[1784] = 1'd0;
    assign memhint[1785] = 1'd0;
    assign memhint[1786] = 1'd0;
    assign memhint[1787] = 1'd0;
    assign memhint[1788] = 1'd0;
    assign memhint[1789] = 1'd0;
    assign memhint[1790] = 1'd0;
    assign memhint[1791] = 1'd0;
    assign memhint[1792] = 1'd0;
    assign memhint[1793] = 1'd0;
    assign memhint[1794] = 1'd1;
    assign memhint[1795] = 1'd1;
    assign memhint[1796] = 1'd0;
    assign memhint[1797] = 1'd0;
    assign memhint[1798] = 1'd0;
    assign memhint[1799] = 1'd0;
    assign memhint[1800] = 1'd0;
    assign memhint[1801] = 1'd0;
    assign memhint[1802] = 1'd0;
    assign memhint[1803] = 1'd0;
    assign memhint[1804] = 1'd0;
    assign memhint[1805] = 1'd0;
    assign memhint[1806] = 1'd1;
    assign memhint[1807] = 1'd1;
    assign memhint[1808] = 1'd0;
    assign memhint[1809] = 1'd0;
    assign memhint[1810] = 1'd0;
    assign memhint[1811] = 1'd0;
    assign memhint[1812] = 1'd0;
    assign memhint[1813] = 1'd1;
    assign memhint[1814] = 1'd1;
    assign memhint[1815] = 1'd0;
    assign memhint[1816] = 1'd0;
    assign memhint[1817] = 1'd0;
    assign memhint[1818] = 1'd0;
    assign memhint[1819] = 1'd0;
    assign memhint[1820] = 1'd0;
    assign memhint[1821] = 1'd0;
    assign memhint[1822] = 1'd0;
    assign memhint[1823] = 1'd0;
    assign memhint[1824] = 1'd0;
    assign memhint[1825] = 1'd0;
    assign memhint[1826] = 1'd0;
    assign memhint[1827] = 1'd0;
    assign memhint[1828] = 1'd0;
    assign memhint[1829] = 1'd0;
    assign memhint[1830] = 1'd0;
    assign memhint[1831] = 1'd0;
    assign memhint[1832] = 1'd0;
    assign memhint[1833] = 1'd0;
    assign memhint[1834] = 1'd1;
    assign memhint[1835] = 1'd1;
    assign memhint[1836] = 1'd0;
    assign memhint[1837] = 1'd1;
    assign memhint[1838] = 1'd1;
    assign memhint[1839] = 1'd0;
    assign memhint[1840] = 1'd0;
    assign memhint[1841] = 1'd0;
    assign memhint[1842] = 1'd0;
    assign memhint[1843] = 1'd0;
    assign memhint[1844] = 1'd0;
    assign memhint[1845] = 1'd0;
    assign memhint[1846] = 1'd0;
    assign memhint[1847] = 1'd0;
    assign memhint[1848] = 1'd0;
    assign memhint[1849] = 1'd0;
    assign memhint[1850] = 1'd0;
    assign memhint[1851] = 1'd0;
    assign memhint[1852] = 1'd1;
    assign memhint[1853] = 1'd1;
    assign memhint[1854] = 1'd0;
    assign memhint[1855] = 1'd0;
    assign memhint[1856] = 1'd0;
    assign memhint[1857] = 1'd0;
    assign memhint[1858] = 1'd0;
    assign memhint[1859] = 1'd0;
    assign memhint[1860] = 1'd1;
    assign memhint[1861] = 1'd1;
    assign memhint[1862] = 1'd0;
    assign memhint[1863] = 1'd0;
    assign memhint[1864] = 1'd0;
    assign memhint[1865] = 1'd0;
    assign memhint[1866] = 1'd1;
    assign memhint[1867] = 1'd1;
    assign memhint[1868] = 1'd0;
    assign memhint[1869] = 1'd0;
    assign memhint[1870] = 1'd0;
    assign memhint[1871] = 1'd0;
    assign memhint[1872] = 1'd0;
    assign memhint[1873] = 1'd0;
    assign memhint[1874] = 1'd0;
    assign memhint[1875] = 1'd0;
    assign memhint[1876] = 1'd0;
    assign memhint[1877] = 1'd0;
    assign memhint[1878] = 1'd0;
    assign memhint[1879] = 1'd0;
    assign memhint[1880] = 1'd0;
    assign memhint[1881] = 1'd0;
    assign memhint[1882] = 1'd0;
    assign memhint[1883] = 1'd1;
    assign memhint[1884] = 1'd1;
    assign memhint[1885] = 1'd0;
    assign memhint[1886] = 1'd0;
    assign memhint[1887] = 1'd0;
    assign memhint[1888] = 1'd0;
    assign memhint[1889] = 1'd0;
    assign memhint[1890] = 1'd0;
    assign memhint[1891] = 1'd0;
    assign memhint[1892] = 1'd0;
    assign memhint[1893] = 1'd0;
    assign memhint[1894] = 1'd0;
    assign memhint[1895] = 1'd0;
    assign memhint[1896] = 1'd0;
    assign memhint[1897] = 1'd0;
    assign memhint[1898] = 1'd0;
    assign memhint[1899] = 1'd0;
    assign memhint[1900] = 1'd1;
    assign memhint[1901] = 1'd1;
    assign memhint[1902] = 1'd0;
    assign memhint[1903] = 1'd0;
    assign memhint[1904] = 1'd0;
    assign memhint[1905] = 1'd0;
    assign memhint[1906] = 1'd0;
    assign memhint[1907] = 1'd0;
    assign memhint[1908] = 1'd0;
    assign memhint[1909] = 1'd0;
    assign memhint[1910] = 1'd0;
    assign memhint[1911] = 1'd0;
    assign memhint[1912] = 1'd0;
    assign memhint[1913] = 1'd0;
    assign memhint[1914] = 1'd0;
    assign memhint[1915] = 1'd1;
    assign memhint[1916] = 1'd1;
    assign memhint[1917] = 1'd0;
    assign memhint[1918] = 1'd0;
    assign memhint[1919] = 1'd0;
    assign memhint[1920] = 1'd0;
    assign memhint[1921] = 1'd0;
    assign memhint[1922] = 1'd0;
    assign memhint[1923] = 1'd0;
    assign memhint[1924] = 1'd0;
    assign memhint[1925] = 1'd0;
    assign memhint[1926] = 1'd0;
    assign memhint[1927] = 1'd0;
    assign memhint[1928] = 1'd0;
    assign memhint[1929] = 1'd0;
    assign memhint[1930] = 1'd0;
    assign memhint[1931] = 1'd0;
    assign memhint[1932] = 1'd0;
    assign memhint[1933] = 1'd1;
    assign memhint[1934] = 1'd1;
    assign memhint[1935] = 1'd0;
    assign memhint[1936] = 1'd0;
    assign memhint[1937] = 1'd0;
    assign memhint[1938] = 1'd0;
    assign memhint[1939] = 1'd0;
    assign memhint[1940] = 1'd0;
    assign memhint[1941] = 1'd0;
    assign memhint[1942] = 1'd0;
    assign memhint[1943] = 1'd0;
    assign memhint[1944] = 1'd0;
    assign memhint[1945] = 1'd0;
    assign memhint[1946] = 1'd0;
    assign memhint[1947] = 1'd0;
    assign memhint[1948] = 1'd0;
    assign memhint[1949] = 1'd0;
    assign memhint[1950] = 1'd0;
    assign memhint[1951] = 1'd1;
    assign memhint[1952] = 1'd0;
    assign memhint[1953] = 1'd0;
    assign memhint[1954] = 1'd0;
    assign memhint[1955] = 1'd0;
    assign memhint[1956] = 1'd0;
    assign memhint[1957] = 1'd0;
    assign memhint[1958] = 1'd0;
    assign memhint[1959] = 1'd0;
    assign memhint[1960] = 1'd1;
    assign memhint[1961] = 1'd1;
    assign memhint[1962] = 1'd0;
    assign memhint[1963] = 1'd0;
    assign memhint[1964] = 1'd0;
    assign memhint[1965] = 1'd0;
    assign memhint[1966] = 1'd0;
    assign memhint[1967] = 1'd0;
    assign memhint[1968] = 1'd0;
    assign memhint[1969] = 1'd0;
    assign memhint[1970] = 1'd0;
    assign memhint[1971] = 1'd0;
    assign memhint[1972] = 1'd0;
    assign memhint[1973] = 1'd0;
    assign memhint[1974] = 1'd0;
    assign memhint[1975] = 1'd0;
    assign memhint[1976] = 1'd0;
    assign memhint[1977] = 1'd0;
    assign memhint[1978] = 1'd0;
    assign memhint[1979] = 1'd0;
    assign memhint[1980] = 1'd0;
    assign memhint[1981] = 1'd0;
    assign memhint[1982] = 1'd0;
    assign memhint[1983] = 1'd0;
    assign memhint[1984] = 1'd0;
    assign memhint[1985] = 1'd0;
    assign memhint[1986] = 1'd1;
    assign memhint[1987] = 1'd1;
    assign memhint[1988] = 1'd0;
    assign memhint[1989] = 1'd1;
    assign memhint[1990] = 1'd1;
    assign memhint[1991] = 1'd0;
    assign memhint[1992] = 1'd0;
    assign memhint[1993] = 1'd0;
    assign memhint[1994] = 1'd0;
    assign memhint[1995] = 1'd0;
    assign memhint[1996] = 1'd0;
    assign memhint[1997] = 1'd0;
    assign memhint[1998] = 1'd0;
    assign memhint[1999] = 1'd0;
    assign memhint[2000] = 1'd0;
    assign memhint[2001] = 1'd0;
    assign memhint[2002] = 1'd0;
    assign memhint[2003] = 1'd0;
    assign memhint[2004] = 1'd0;
    assign memhint[2005] = 1'd0;
    assign memhint[2006] = 1'd0;
    assign memhint[2007] = 1'd0;
    assign memhint[2008] = 1'd0;
    assign memhint[2009] = 1'd0;
    assign memhint[2010] = 1'd0;
    assign memhint[2011] = 1'd1;
    assign memhint[2012] = 1'd1;
    assign memhint[2013] = 1'd0;
    assign memhint[2014] = 1'd0;
    assign memhint[2015] = 1'd0;
    assign memhint[2016] = 1'd0;
    assign memhint[2017] = 1'd0;
    assign memhint[2018] = 1'd0;
    assign memhint[2019] = 1'd0;
    assign memhint[2020] = 1'd0;
    assign memhint[2021] = 1'd0;
    assign memhint[2022] = 1'd0;
    assign memhint[2023] = 1'd0;
    assign memhint[2024] = 1'd0;
    assign memhint[2025] = 1'd0;
    assign memhint[2026] = 1'd0;
    assign memhint[2027] = 1'd0;
    assign memhint[2028] = 1'd0;
    assign memhint[2029] = 1'd1;
    assign memhint[2030] = 1'd1;
    assign memhint[2031] = 1'd0;
    assign memhint[2032] = 1'd0;
    assign memhint[2033] = 1'd0;
    assign memhint[2034] = 1'd0;
    assign memhint[2035] = 1'd0;
    assign memhint[2036] = 1'd0;
    assign memhint[2037] = 1'd0;
    assign memhint[2038] = 1'd0;
    assign memhint[2039] = 1'd0;
    assign memhint[2040] = 1'd0;
    assign memhint[2041] = 1'd0;
    assign memhint[2042] = 1'd0;
    assign memhint[2043] = 1'd0;
    assign memhint[2044] = 1'd0;
    assign memhint[2045] = 1'd0;
    assign memhint[2046] = 1'd0;
    assign memhint[2047] = 1'd1;
    assign memhint[2048] = 1'd1;
    assign memhint[2049] = 1'd0;
    assign memhint[2050] = 1'd0;
    assign memhint[2051] = 1'd0;
    assign memhint[2052] = 1'd0;
    assign memhint[2053] = 1'd0;
    assign memhint[2054] = 1'd0;
    assign memhint[2055] = 1'd0;
    assign memhint[2056] = 1'd1;
    assign memhint[2057] = 1'd1;
    assign memhint[2058] = 1'd0;
    assign memhint[2059] = 1'd1;
    assign memhint[2060] = 1'd1;
    assign memhint[2061] = 1'd0;
    assign memhint[2062] = 1'd0;
    assign memhint[2063] = 1'd0;
    assign memhint[2064] = 1'd0;
    assign memhint[2065] = 1'd0;
    assign memhint[2066] = 1'd0;
    assign memhint[2067] = 1'd0;
    assign memhint[2068] = 1'd0;
    assign memhint[2069] = 1'd0;
    assign memhint[2070] = 1'd0;
    assign memhint[2071] = 1'd0;
    assign memhint[2072] = 1'd1;
    assign memhint[2073] = 1'd1;
    assign memhint[2074] = 1'd0;
    assign memhint[2075] = 1'd0;
    assign memhint[2076] = 1'd0;
    assign memhint[2077] = 1'd0;
    assign memhint[2078] = 1'd0;
    assign memhint[2079] = 1'd0;
    assign memhint[2080] = 1'd0;
    assign memhint[2081] = 1'd1;
    assign memhint[2082] = 1'd1;
    assign memhint[2083] = 1'd0;
    assign memhint[2084] = 1'd0;
    assign memhint[2085] = 1'd0;
    assign memhint[2086] = 1'd0;
    assign memhint[2087] = 1'd0;
    assign memhint[2088] = 1'd0;
    assign memhint[2089] = 1'd0;
    assign memhint[2090] = 1'd0;
    assign memhint[2091] = 1'd0;
    assign memhint[2092] = 1'd0;
    assign memhint[2093] = 1'd0;
    assign memhint[2094] = 1'd0;
    assign memhint[2095] = 1'd0;
    assign memhint[2096] = 1'd0;
    assign memhint[2097] = 1'd0;
    assign memhint[2098] = 1'd0;
    assign memhint[2099] = 1'd0;
    assign memhint[2100] = 1'd1;
    assign memhint[2101] = 1'd0;
    assign memhint[2102] = 1'd0;
    assign memhint[2103] = 1'd0;
    assign memhint[2104] = 1'd0;
    assign memhint[2105] = 1'd0;
    assign memhint[2106] = 1'd0;
    assign memhint[2107] = 1'd0;
    assign memhint[2108] = 1'd0;
    assign memhint[2109] = 1'd0;
    assign memhint[2110] = 1'd0;
    assign memhint[2111] = 1'd0;
    assign memhint[2112] = 1'd0;
    assign memhint[2113] = 1'd0;
    assign memhint[2114] = 1'd0;
    assign memhint[2115] = 1'd0;
    assign memhint[2116] = 1'd0;
    assign memhint[2117] = 1'd0;
    assign memhint[2118] = 1'd0;
    assign memhint[2119] = 1'd1;
    assign memhint[2120] = 1'd1;
    assign memhint[2121] = 1'd0;
    assign memhint[2122] = 1'd0;
    assign memhint[2123] = 1'd0;
    assign memhint[2124] = 1'd0;
    assign memhint[2125] = 1'd0;
    assign memhint[2126] = 1'd0;
    assign memhint[2127] = 1'd0;
    assign memhint[2128] = 1'd0;
    assign memhint[2129] = 1'd0;
    assign memhint[2130] = 1'd0;
    assign memhint[2131] = 1'd1;
    assign memhint[2132] = 1'd1;
    assign memhint[2133] = 1'd0;
    assign memhint[2134] = 1'd0;
    assign memhint[2135] = 1'd0;
    assign memhint[2136] = 1'd0;
    assign memhint[2137] = 1'd0;
    assign memhint[2138] = 1'd0;
    assign memhint[2139] = 1'd0;
    assign memhint[2140] = 1'd0;
    assign memhint[2141] = 1'd0;
    assign memhint[2142] = 1'd0;
    assign memhint[2143] = 1'd0;
    assign memhint[2144] = 1'd0;
    assign memhint[2145] = 1'd0;
    assign memhint[2146] = 1'd0;
    assign memhint[2147] = 1'd0;
    assign memhint[2148] = 1'd0;
    assign memhint[2149] = 1'd1;
    assign memhint[2150] = 1'd1;
    assign memhint[2151] = 1'd0;
    assign memhint[2152] = 1'd0;
    assign memhint[2153] = 1'd0;
    assign memhint[2154] = 1'd0;
    assign memhint[2155] = 1'd0;
    assign memhint[2156] = 1'd0;
    assign memhint[2157] = 1'd0;
    assign memhint[2158] = 1'd0;
    assign memhint[2159] = 1'd0;
    assign memhint[2160] = 1'd0;
    assign memhint[2161] = 1'd0;
    assign memhint[2162] = 1'd0;
    assign memhint[2163] = 1'd0;
    assign memhint[2164] = 1'd0;
    assign memhint[2165] = 1'd0;
    assign memhint[2166] = 1'd0;
    assign memhint[2167] = 1'd1;
    assign memhint[2168] = 1'd1;
    assign memhint[2169] = 1'd0;
    assign memhint[2170] = 1'd0;
    assign memhint[2171] = 1'd0;
    assign memhint[2172] = 1'd0;
    assign memhint[2173] = 1'd0;
    assign memhint[2174] = 1'd0;
    assign memhint[2175] = 1'd0;
    assign memhint[2176] = 1'd0;
    assign memhint[2177] = 1'd0;
    assign memhint[2178] = 1'd0;
    assign memhint[2179] = 1'd1;
    assign memhint[2180] = 1'd1;
    assign memhint[2181] = 1'd0;
    assign memhint[2182] = 1'd0;
    assign memhint[2183] = 1'd0;
    assign memhint[2184] = 1'd0;
    assign memhint[2185] = 1'd0;
    assign memhint[2186] = 1'd1;
    assign memhint[2187] = 1'd1;
    assign memhint[2188] = 1'd0;
    assign memhint[2189] = 1'd0;
    assign memhint[2190] = 1'd0;
    assign memhint[2191] = 1'd0;
    assign memhint[2192] = 1'd0;
    assign memhint[2193] = 1'd0;
    assign memhint[2194] = 1'd0;
    assign memhint[2195] = 1'd0;
    assign memhint[2196] = 1'd0;
    assign memhint[2197] = 1'd0;
    assign memhint[2198] = 1'd0;
    assign memhint[2199] = 1'd0;
    assign memhint[2200] = 1'd0;
    assign memhint[2201] = 1'd0;
    assign memhint[2202] = 1'd0;
    assign memhint[2203] = 1'd0;
    assign memhint[2204] = 1'd0;
    assign memhint[2205] = 1'd0;
    assign memhint[2206] = 1'd0;
    assign memhint[2207] = 1'd1;
    assign memhint[2208] = 1'd1;
    assign memhint[2209] = 1'd0;
    assign memhint[2210] = 1'd1;
    assign memhint[2211] = 1'd1;
    assign memhint[2212] = 1'd0;
    assign memhint[2213] = 1'd0;
    assign memhint[2214] = 1'd0;
    assign memhint[2215] = 1'd0;
    assign memhint[2216] = 1'd0;
    assign memhint[2217] = 1'd0;
    assign memhint[2218] = 1'd0;
    assign memhint[2219] = 1'd0;
    assign memhint[2220] = 1'd0;
    assign memhint[2221] = 1'd0;
    assign memhint[2222] = 1'd0;
    assign memhint[2223] = 1'd0;
    assign memhint[2224] = 1'd0;
    assign memhint[2225] = 1'd1;
    assign memhint[2226] = 1'd1;
    assign memhint[2227] = 1'd0;
    assign memhint[2228] = 1'd0;
    assign memhint[2229] = 1'd0;
    assign memhint[2230] = 1'd0;
    assign memhint[2231] = 1'd0;
    assign memhint[2232] = 1'd0;
    assign memhint[2233] = 1'd1;
    assign memhint[2234] = 1'd1;
    assign memhint[2235] = 1'd0;
    assign memhint[2236] = 1'd0;
    assign memhint[2237] = 1'd0;
    assign memhint[2238] = 1'd0;
    assign memhint[2239] = 1'd1;
    assign memhint[2240] = 1'd1;
    assign memhint[2241] = 1'd0;
    assign memhint[2242] = 1'd0;
    assign memhint[2243] = 1'd0;
    assign memhint[2244] = 1'd0;
    assign memhint[2245] = 1'd0;
    assign memhint[2246] = 1'd0;
    assign memhint[2247] = 1'd0;
    assign memhint[2248] = 1'd0;
    assign memhint[2249] = 1'd0;
    assign memhint[2250] = 1'd0;
    assign memhint[2251] = 1'd0;
    assign memhint[2252] = 1'd0;
    assign memhint[2253] = 1'd0;
    assign memhint[2254] = 1'd0;
    assign memhint[2255] = 1'd0;
    assign memhint[2256] = 1'd1;
    assign memhint[2257] = 1'd1;
    assign memhint[2258] = 1'd0;
    assign memhint[2259] = 1'd0;
    assign memhint[2260] = 1'd0;
    assign memhint[2261] = 1'd0;
    assign memhint[2262] = 1'd0;
    assign memhint[2263] = 1'd0;
    assign memhint[2264] = 1'd0;
    assign memhint[2265] = 1'd0;
    assign memhint[2266] = 1'd0;
    assign memhint[2267] = 1'd0;
    assign memhint[2268] = 1'd0;
    assign memhint[2269] = 1'd0;
    assign memhint[2270] = 1'd0;
    assign memhint[2271] = 1'd0;
    assign memhint[2272] = 1'd0;
    assign memhint[2273] = 1'd1;
    assign memhint[2274] = 1'd1;
    assign memhint[2275] = 1'd0;
    assign memhint[2276] = 1'd0;
    assign memhint[2277] = 1'd0;
    assign memhint[2278] = 1'd0;
    assign memhint[2279] = 1'd0;
    assign memhint[2280] = 1'd0;
    assign memhint[2281] = 1'd0;
    assign memhint[2282] = 1'd0;
    assign memhint[2283] = 1'd0;
    assign memhint[2284] = 1'd0;
    assign memhint[2285] = 1'd0;
    assign memhint[2286] = 1'd0;
    assign memhint[2287] = 1'd0;
    assign memhint[2288] = 1'd1;
    assign memhint[2289] = 1'd1;
    assign memhint[2290] = 1'd0;
    assign memhint[2291] = 1'd0;
    assign memhint[2292] = 1'd0;
    assign memhint[2293] = 1'd0;
    assign memhint[2294] = 1'd0;
    assign memhint[2295] = 1'd0;
    assign memhint[2296] = 1'd0;
    assign memhint[2297] = 1'd0;
    assign memhint[2298] = 1'd0;
    assign memhint[2299] = 1'd0;
    assign memhint[2300] = 1'd0;
    assign memhint[2301] = 1'd0;
    assign memhint[2302] = 1'd0;
    assign memhint[2303] = 1'd0;
    assign memhint[2304] = 1'd0;
    assign memhint[2305] = 1'd1;
    assign memhint[2306] = 1'd1;
    assign memhint[2307] = 1'd0;
    assign memhint[2308] = 1'd0;
    assign memhint[2309] = 1'd0;
    assign memhint[2310] = 1'd0;
    assign memhint[2311] = 1'd0;
    assign memhint[2312] = 1'd0;
    assign memhint[2313] = 1'd0;
    assign memhint[2314] = 1'd0;
    assign memhint[2315] = 1'd0;
    assign memhint[2316] = 1'd0;
    assign memhint[2317] = 1'd0;
    assign memhint[2318] = 1'd0;
    assign memhint[2319] = 1'd0;
    assign memhint[2320] = 1'd0;
    assign memhint[2321] = 1'd0;
    assign memhint[2322] = 1'd0;
    assign memhint[2323] = 1'd0;
    assign memhint[2324] = 1'd0;
    assign memhint[2325] = 1'd0;
    assign memhint[2326] = 1'd0;
    assign memhint[2327] = 1'd0;
    assign memhint[2328] = 1'd0;
    assign memhint[2329] = 1'd0;
    assign memhint[2330] = 1'd0;
    assign memhint[2331] = 1'd0;
    assign memhint[2332] = 1'd0;
    assign memhint[2333] = 1'd1;
    assign memhint[2334] = 1'd1;
    assign memhint[2335] = 1'd0;
    assign memhint[2336] = 1'd0;
    assign memhint[2337] = 1'd0;
    assign memhint[2338] = 1'd0;
    assign memhint[2339] = 1'd0;
    assign memhint[2340] = 1'd0;
    assign memhint[2341] = 1'd0;
    assign memhint[2342] = 1'd0;
    assign memhint[2343] = 1'd0;
    assign memhint[2344] = 1'd0;
    assign memhint[2345] = 1'd0;
    assign memhint[2346] = 1'd0;
    assign memhint[2347] = 1'd0;
    assign memhint[2348] = 1'd0;
    assign memhint[2349] = 1'd0;
    assign memhint[2350] = 1'd0;
    assign memhint[2351] = 1'd0;
    assign memhint[2352] = 1'd0;
    assign memhint[2353] = 1'd0;
    assign memhint[2354] = 1'd0;
    assign memhint[2355] = 1'd0;
    assign memhint[2356] = 1'd0;
    assign memhint[2357] = 1'd0;
    assign memhint[2358] = 1'd1;
    assign memhint[2359] = 1'd1;
    assign memhint[2360] = 1'd0;
    assign memhint[2361] = 1'd0;
    assign memhint[2362] = 1'd0;
    assign memhint[2363] = 1'd1;
    assign memhint[2364] = 1'd1;
    assign memhint[2365] = 1'd0;
    assign memhint[2366] = 1'd0;
    assign memhint[2367] = 1'd0;
    assign memhint[2368] = 1'd0;
    assign memhint[2369] = 1'd0;
    assign memhint[2370] = 1'd0;
    assign memhint[2371] = 1'd0;
    assign memhint[2372] = 1'd0;
    assign memhint[2373] = 1'd0;
    assign memhint[2374] = 1'd0;
    assign memhint[2375] = 1'd0;
    assign memhint[2376] = 1'd0;
    assign memhint[2377] = 1'd0;
    assign memhint[2378] = 1'd0;
    assign memhint[2379] = 1'd0;
    assign memhint[2380] = 1'd0;
    assign memhint[2381] = 1'd0;
    assign memhint[2382] = 1'd0;
    assign memhint[2383] = 1'd0;
    assign memhint[2384] = 1'd1;
    assign memhint[2385] = 1'd1;
    assign memhint[2386] = 1'd0;
    assign memhint[2387] = 1'd0;
    assign memhint[2388] = 1'd0;
    assign memhint[2389] = 1'd0;
    assign memhint[2390] = 1'd0;
    assign memhint[2391] = 1'd0;
    assign memhint[2392] = 1'd0;
    assign memhint[2393] = 1'd0;
    assign memhint[2394] = 1'd0;
    assign memhint[2395] = 1'd0;
    assign memhint[2396] = 1'd0;
    assign memhint[2397] = 1'd0;
    assign memhint[2398] = 1'd0;
    assign memhint[2399] = 1'd0;
    assign memhint[2400] = 1'd0;
    assign memhint[2401] = 1'd1;
    assign memhint[2402] = 1'd1;
    assign memhint[2403] = 1'd0;
    assign memhint[2404] = 1'd0;
    assign memhint[2405] = 1'd0;
    assign memhint[2406] = 1'd0;
    assign memhint[2407] = 1'd0;
    assign memhint[2408] = 1'd0;
    assign memhint[2409] = 1'd0;
    assign memhint[2410] = 1'd0;
    assign memhint[2411] = 1'd0;
    assign memhint[2412] = 1'd0;
    assign memhint[2413] = 1'd0;
    assign memhint[2414] = 1'd0;
    assign memhint[2415] = 1'd0;
    assign memhint[2416] = 1'd0;
    assign memhint[2417] = 1'd0;
    assign memhint[2418] = 1'd0;
    assign memhint[2419] = 1'd0;
    assign memhint[2420] = 1'd0;
    assign memhint[2421] = 1'd1;
    assign memhint[2422] = 1'd1;
    assign memhint[2423] = 1'd0;
    assign memhint[2424] = 1'd0;
    assign memhint[2425] = 1'd0;
    assign memhint[2426] = 1'd0;
    assign memhint[2427] = 1'd0;
    assign memhint[2428] = 1'd0;
    assign memhint[2429] = 1'd1;
    assign memhint[2430] = 1'd1;
    assign memhint[2431] = 1'd0;
    assign memhint[2432] = 1'd0;
    assign memhint[2433] = 1'd1;
    assign memhint[2434] = 1'd1;
    assign memhint[2435] = 1'd0;
    assign memhint[2436] = 1'd0;
    assign memhint[2437] = 1'd0;
    assign memhint[2438] = 1'd0;
    assign memhint[2439] = 1'd0;
    assign memhint[2440] = 1'd0;
    assign memhint[2441] = 1'd0;
    assign memhint[2442] = 1'd0;
    assign memhint[2443] = 1'd0;
    assign memhint[2444] = 1'd0;
    assign memhint[2445] = 1'd1;
    assign memhint[2446] = 1'd1;
    assign memhint[2447] = 1'd0;
    assign memhint[2448] = 1'd0;
    assign memhint[2449] = 1'd0;
    assign memhint[2450] = 1'd0;
    assign memhint[2451] = 1'd0;
    assign memhint[2452] = 1'd0;
    assign memhint[2453] = 1'd1;
    assign memhint[2454] = 1'd1;
    assign memhint[2455] = 1'd1;
    assign memhint[2456] = 1'd0;
    assign memhint[2457] = 1'd0;
    assign memhint[2458] = 1'd0;
    assign memhint[2459] = 1'd0;
    assign memhint[2460] = 1'd0;
    assign memhint[2461] = 1'd0;
    assign memhint[2462] = 1'd0;
    assign memhint[2463] = 1'd0;
    assign memhint[2464] = 1'd0;
    assign memhint[2465] = 1'd0;
    assign memhint[2466] = 1'd0;
    assign memhint[2467] = 1'd0;
    assign memhint[2468] = 1'd0;
    assign memhint[2469] = 1'd0;
    assign memhint[2470] = 1'd0;
    assign memhint[2471] = 1'd0;
    assign memhint[2472] = 1'd0;
    assign memhint[2473] = 1'd0;
    assign memhint[2474] = 1'd0;
    assign memhint[2475] = 1'd0;
    assign memhint[2476] = 1'd0;
    assign memhint[2477] = 1'd0;
    assign memhint[2478] = 1'd0;
    assign memhint[2479] = 1'd0;
    assign memhint[2480] = 1'd0;
    assign memhint[2481] = 1'd0;
    assign memhint[2482] = 1'd0;
    assign memhint[2483] = 1'd0;
    assign memhint[2484] = 1'd0;
    assign memhint[2485] = 1'd0;
    assign memhint[2486] = 1'd0;
    assign memhint[2487] = 1'd0;
    assign memhint[2488] = 1'd0;
    assign memhint[2489] = 1'd0;
    assign memhint[2490] = 1'd0;
    assign memhint[2491] = 1'd0;
    assign memhint[2492] = 1'd1;
    assign memhint[2493] = 1'd1;
    assign memhint[2494] = 1'd0;
    assign memhint[2495] = 1'd0;
    assign memhint[2496] = 1'd0;
    assign memhint[2497] = 1'd0;
    assign memhint[2498] = 1'd0;
    assign memhint[2499] = 1'd0;
    assign memhint[2500] = 1'd0;
    assign memhint[2501] = 1'd0;
    assign memhint[2502] = 1'd0;
    assign memhint[2503] = 1'd1;
    assign memhint[2504] = 1'd1;
    assign memhint[2505] = 1'd0;
    assign memhint[2506] = 1'd0;
    assign memhint[2507] = 1'd0;
    assign memhint[2508] = 1'd0;
    assign memhint[2509] = 1'd0;
    assign memhint[2510] = 1'd0;
    assign memhint[2511] = 1'd0;
    assign memhint[2512] = 1'd0;
    assign memhint[2513] = 1'd0;
    assign memhint[2514] = 1'd0;
    assign memhint[2515] = 1'd0;
    assign memhint[2516] = 1'd0;
    assign memhint[2517] = 1'd0;
    assign memhint[2518] = 1'd0;
    assign memhint[2519] = 1'd0;
    assign memhint[2520] = 1'd0;
    assign memhint[2521] = 1'd0;
    assign memhint[2522] = 1'd0;
    assign memhint[2523] = 1'd1;
    assign memhint[2524] = 1'd1;
    assign memhint[2525] = 1'd0;
    assign memhint[2526] = 1'd0;
    assign memhint[2527] = 1'd0;
    assign memhint[2528] = 1'd0;
    assign memhint[2529] = 1'd0;
    assign memhint[2530] = 1'd0;
    assign memhint[2531] = 1'd0;
    assign memhint[2532] = 1'd0;
    assign memhint[2533] = 1'd0;
    assign memhint[2534] = 1'd0;
    assign memhint[2535] = 1'd0;
    assign memhint[2536] = 1'd0;
    assign memhint[2537] = 1'd0;
    assign memhint[2538] = 1'd0;
    assign memhint[2539] = 1'd0;
    assign memhint[2540] = 1'd1;
    assign memhint[2541] = 1'd1;
    assign memhint[2542] = 1'd0;
    assign memhint[2543] = 1'd0;
    assign memhint[2544] = 1'd0;
    assign memhint[2545] = 1'd0;
    assign memhint[2546] = 1'd0;
    assign memhint[2547] = 1'd0;
    assign memhint[2548] = 1'd0;
    assign memhint[2549] = 1'd0;
    assign memhint[2550] = 1'd0;
    assign memhint[2551] = 1'd0;
    assign memhint[2552] = 1'd1;
    assign memhint[2553] = 1'd1;
    assign memhint[2554] = 1'd0;
    assign memhint[2555] = 1'd0;
    assign memhint[2556] = 1'd0;
    assign memhint[2557] = 1'd0;
    assign memhint[2558] = 1'd0;
    assign memhint[2559] = 1'd1;
    assign memhint[2560] = 1'd1;
    assign memhint[2561] = 1'd0;
    assign memhint[2562] = 1'd0;
    assign memhint[2563] = 1'd0;
    assign memhint[2564] = 1'd0;
    assign memhint[2565] = 1'd0;
    assign memhint[2566] = 1'd0;
    assign memhint[2567] = 1'd0;
    assign memhint[2568] = 1'd0;
    assign memhint[2569] = 1'd0;
    assign memhint[2570] = 1'd0;
    assign memhint[2571] = 1'd0;
    assign memhint[2572] = 1'd0;
    assign memhint[2573] = 1'd0;
    assign memhint[2574] = 1'd0;
    assign memhint[2575] = 1'd0;
    assign memhint[2576] = 1'd0;
    assign memhint[2577] = 1'd0;
    assign memhint[2578] = 1'd0;
    assign memhint[2579] = 1'd1;
    assign memhint[2580] = 1'd1;
    assign memhint[2581] = 1'd0;
    assign memhint[2582] = 1'd0;
    assign memhint[2583] = 1'd0;
    assign memhint[2584] = 1'd1;
    assign memhint[2585] = 1'd1;
    assign memhint[2586] = 1'd0;
    assign memhint[2587] = 1'd0;
    assign memhint[2588] = 1'd0;
    assign memhint[2589] = 1'd0;
    assign memhint[2590] = 1'd0;
    assign memhint[2591] = 1'd0;
    assign memhint[2592] = 1'd0;
    assign memhint[2593] = 1'd0;
    assign memhint[2594] = 1'd0;
    assign memhint[2595] = 1'd0;
    assign memhint[2596] = 1'd0;
    assign memhint[2597] = 1'd0;
    assign memhint[2598] = 1'd0;
    assign memhint[2599] = 1'd1;
    assign memhint[2600] = 1'd1;
    assign memhint[2601] = 1'd0;
    assign memhint[2602] = 1'd0;
    assign memhint[2603] = 1'd0;
    assign memhint[2604] = 1'd0;
    assign memhint[2605] = 1'd1;
    assign memhint[2606] = 1'd1;
    assign memhint[2607] = 1'd0;
    assign memhint[2608] = 1'd0;
    assign memhint[2609] = 1'd0;
    assign memhint[2610] = 1'd0;
    assign memhint[2611] = 1'd0;
    assign memhint[2612] = 1'd0;
    assign memhint[2613] = 1'd1;
    assign memhint[2614] = 1'd1;
    assign memhint[2615] = 1'd0;
    assign memhint[2616] = 1'd0;
    assign memhint[2617] = 1'd0;
    assign memhint[2618] = 1'd0;
    assign memhint[2619] = 1'd0;
    assign memhint[2620] = 1'd0;
    assign memhint[2621] = 1'd0;
    assign memhint[2622] = 1'd0;
    assign memhint[2623] = 1'd0;
    assign memhint[2624] = 1'd0;
    assign memhint[2625] = 1'd0;
    assign memhint[2626] = 1'd0;
    assign memhint[2627] = 1'd0;
    assign memhint[2628] = 1'd0;
    assign memhint[2629] = 1'd1;
    assign memhint[2630] = 1'd1;
    assign memhint[2631] = 1'd0;
    assign memhint[2632] = 1'd0;
    assign memhint[2633] = 1'd0;
    assign memhint[2634] = 1'd0;
    assign memhint[2635] = 1'd0;
    assign memhint[2636] = 1'd0;
    assign memhint[2637] = 1'd0;
    assign memhint[2638] = 1'd0;
    assign memhint[2639] = 1'd0;
    assign memhint[2640] = 1'd0;
    assign memhint[2641] = 1'd0;
    assign memhint[2642] = 1'd0;
    assign memhint[2643] = 1'd0;
    assign memhint[2644] = 1'd0;
    assign memhint[2645] = 1'd0;
    assign memhint[2646] = 1'd1;
    assign memhint[2647] = 1'd1;
    assign memhint[2648] = 1'd0;
    assign memhint[2649] = 1'd0;
    assign memhint[2650] = 1'd0;
    assign memhint[2651] = 1'd0;
    assign memhint[2652] = 1'd0;
    assign memhint[2653] = 1'd0;
    assign memhint[2654] = 1'd0;
    assign memhint[2655] = 1'd0;
    assign memhint[2656] = 1'd0;
    assign memhint[2657] = 1'd0;
    assign memhint[2658] = 1'd0;
    assign memhint[2659] = 1'd0;
    assign memhint[2660] = 1'd0;
    assign memhint[2661] = 1'd1;
    assign memhint[2662] = 1'd1;
    assign memhint[2663] = 1'd0;
    assign memhint[2664] = 1'd0;
    assign memhint[2665] = 1'd0;
    assign memhint[2666] = 1'd0;
    assign memhint[2667] = 1'd0;
    assign memhint[2668] = 1'd0;
    assign memhint[2669] = 1'd0;
    assign memhint[2670] = 1'd0;
    assign memhint[2671] = 1'd0;
    assign memhint[2672] = 1'd0;
    assign memhint[2673] = 1'd0;
    assign memhint[2674] = 1'd0;
    assign memhint[2675] = 1'd0;
    assign memhint[2676] = 1'd0;
    assign memhint[2677] = 1'd0;
    assign memhint[2678] = 1'd1;
    assign memhint[2679] = 1'd1;
    assign memhint[2680] = 1'd0;
    assign memhint[2681] = 1'd0;
    assign memhint[2682] = 1'd0;
    assign memhint[2683] = 1'd0;
    assign memhint[2684] = 1'd0;
    assign memhint[2685] = 1'd0;
    assign memhint[2686] = 1'd0;
    assign memhint[2687] = 1'd0;
    assign memhint[2688] = 1'd0;
    assign memhint[2689] = 1'd0;
    assign memhint[2690] = 1'd0;
    assign memhint[2691] = 1'd0;
    assign memhint[2692] = 1'd0;
    assign memhint[2693] = 1'd0;
    assign memhint[2694] = 1'd0;
    assign memhint[2695] = 1'd0;
    assign memhint[2696] = 1'd0;
    assign memhint[2697] = 1'd0;
    assign memhint[2698] = 1'd0;
    assign memhint[2699] = 1'd0;
    assign memhint[2700] = 1'd0;
    assign memhint[2701] = 1'd0;
    assign memhint[2702] = 1'd0;
    assign memhint[2703] = 1'd0;
    assign memhint[2704] = 1'd0;
    assign memhint[2705] = 1'd0;
    assign memhint[2706] = 1'd1;
    assign memhint[2707] = 1'd1;
    assign memhint[2708] = 1'd0;
    assign memhint[2709] = 1'd0;
    assign memhint[2710] = 1'd0;
    assign memhint[2711] = 1'd0;
    assign memhint[2712] = 1'd0;
    assign memhint[2713] = 1'd0;
    assign memhint[2714] = 1'd0;
    assign memhint[2715] = 1'd0;
    assign memhint[2716] = 1'd0;
    assign memhint[2717] = 1'd0;
    assign memhint[2718] = 1'd0;
    assign memhint[2719] = 1'd0;
    assign memhint[2720] = 1'd0;
    assign memhint[2721] = 1'd0;
    assign memhint[2722] = 1'd0;
    assign memhint[2723] = 1'd0;
    assign memhint[2724] = 1'd0;
    assign memhint[2725] = 1'd0;
    assign memhint[2726] = 1'd0;
    assign memhint[2727] = 1'd0;
    assign memhint[2728] = 1'd0;
    assign memhint[2729] = 1'd0;
    assign memhint[2730] = 1'd0;
    assign memhint[2731] = 1'd1;
    assign memhint[2732] = 1'd1;
    assign memhint[2733] = 1'd0;
    assign memhint[2734] = 1'd0;
    assign memhint[2735] = 1'd0;
    assign memhint[2736] = 1'd1;
    assign memhint[2737] = 1'd1;
    assign memhint[2738] = 1'd0;
    assign memhint[2739] = 1'd0;
    assign memhint[2740] = 1'd0;
    assign memhint[2741] = 1'd0;
    assign memhint[2742] = 1'd0;
    assign memhint[2743] = 1'd0;
    assign memhint[2744] = 1'd0;
    assign memhint[2745] = 1'd0;
    assign memhint[2746] = 1'd0;
    assign memhint[2747] = 1'd0;
    assign memhint[2748] = 1'd0;
    assign memhint[2749] = 1'd0;
    assign memhint[2750] = 1'd0;
    assign memhint[2751] = 1'd0;
    assign memhint[2752] = 1'd0;
    assign memhint[2753] = 1'd0;
    assign memhint[2754] = 1'd0;
    assign memhint[2755] = 1'd0;
    assign memhint[2756] = 1'd0;
    assign memhint[2757] = 1'd0;
    assign memhint[2758] = 1'd1;
    assign memhint[2759] = 1'd1;
    assign memhint[2760] = 1'd0;
    assign memhint[2761] = 1'd0;
    assign memhint[2762] = 1'd0;
    assign memhint[2763] = 1'd0;
    assign memhint[2764] = 1'd0;
    assign memhint[2765] = 1'd0;
    assign memhint[2766] = 1'd0;
    assign memhint[2767] = 1'd0;
    assign memhint[2768] = 1'd0;
    assign memhint[2769] = 1'd0;
    assign memhint[2770] = 1'd0;
    assign memhint[2771] = 1'd0;
    assign memhint[2772] = 1'd0;
    assign memhint[2773] = 1'd0;
    assign memhint[2774] = 1'd1;
    assign memhint[2775] = 1'd1;
    assign memhint[2776] = 1'd0;
    assign memhint[2777] = 1'd0;
    assign memhint[2778] = 1'd0;
    assign memhint[2779] = 1'd0;
    assign memhint[2780] = 1'd0;
    assign memhint[2781] = 1'd0;
    assign memhint[2782] = 1'd0;
    assign memhint[2783] = 1'd0;
    assign memhint[2784] = 1'd0;
    assign memhint[2785] = 1'd0;
    assign memhint[2786] = 1'd0;
    assign memhint[2787] = 1'd0;
    assign memhint[2788] = 1'd0;
    assign memhint[2789] = 1'd0;
    assign memhint[2790] = 1'd0;
    assign memhint[2791] = 1'd0;
    assign memhint[2792] = 1'd0;
    assign memhint[2793] = 1'd0;
    assign memhint[2794] = 1'd1;
    assign memhint[2795] = 1'd1;
    assign memhint[2796] = 1'd0;
    assign memhint[2797] = 1'd0;
    assign memhint[2798] = 1'd0;
    assign memhint[2799] = 1'd0;
    assign memhint[2800] = 1'd0;
    assign memhint[2801] = 1'd0;
    assign memhint[2802] = 1'd1;
    assign memhint[2803] = 1'd1;
    assign memhint[2804] = 1'd0;
    assign memhint[2805] = 1'd0;
    assign memhint[2806] = 1'd0;
    assign memhint[2807] = 1'd1;
    assign memhint[2808] = 1'd1;
    assign memhint[2809] = 1'd0;
    assign memhint[2810] = 1'd0;
    assign memhint[2811] = 1'd0;
    assign memhint[2812] = 1'd0;
    assign memhint[2813] = 1'd0;
    assign memhint[2814] = 1'd0;
    assign memhint[2815] = 1'd0;
    assign memhint[2816] = 1'd0;
    assign memhint[2817] = 1'd0;
    assign memhint[2818] = 1'd1;
    assign memhint[2819] = 1'd1;
    assign memhint[2820] = 1'd0;
    assign memhint[2821] = 1'd0;
    assign memhint[2822] = 1'd0;
    assign memhint[2823] = 1'd0;
    assign memhint[2824] = 1'd0;
    assign memhint[2825] = 1'd0;
    assign memhint[2826] = 1'd1;
    assign memhint[2827] = 1'd1;
    assign memhint[2828] = 1'd0;
    assign memhint[2829] = 1'd0;
    assign memhint[2830] = 1'd0;
    assign memhint[2831] = 1'd0;
    assign memhint[2832] = 1'd0;
    assign memhint[2833] = 1'd0;
    assign memhint[2834] = 1'd0;
    assign memhint[2835] = 1'd0;
    assign memhint[2836] = 1'd0;
    assign memhint[2837] = 1'd0;
    assign memhint[2838] = 1'd0;
    assign memhint[2839] = 1'd0;
    assign memhint[2840] = 1'd0;
    assign memhint[2841] = 1'd0;
    assign memhint[2842] = 1'd0;
    assign memhint[2843] = 1'd0;
    assign memhint[2844] = 1'd0;
    assign memhint[2845] = 1'd0;
    assign memhint[2846] = 1'd0;
    assign memhint[2847] = 1'd0;
    assign memhint[2848] = 1'd0;
    assign memhint[2849] = 1'd0;
    assign memhint[2850] = 1'd0;
    assign memhint[2851] = 1'd0;
    assign memhint[2852] = 1'd0;
    assign memhint[2853] = 1'd0;
    assign memhint[2854] = 1'd0;
    assign memhint[2855] = 1'd0;
    assign memhint[2856] = 1'd0;
    assign memhint[2857] = 1'd0;
    assign memhint[2858] = 1'd0;
    assign memhint[2859] = 1'd0;
    assign memhint[2860] = 1'd0;
    assign memhint[2861] = 1'd0;
    assign memhint[2862] = 1'd0;
    assign memhint[2863] = 1'd0;
    assign memhint[2864] = 1'd0;
    assign memhint[2865] = 1'd1;
    assign memhint[2866] = 1'd1;
    assign memhint[2867] = 1'd0;
    assign memhint[2868] = 1'd0;
    assign memhint[2869] = 1'd0;
    assign memhint[2870] = 1'd0;
    assign memhint[2871] = 1'd0;
    assign memhint[2872] = 1'd0;
    assign memhint[2873] = 1'd0;
    assign memhint[2874] = 1'd0;
    assign memhint[2875] = 1'd0;
    assign memhint[2876] = 1'd1;
    assign memhint[2877] = 1'd1;
    assign memhint[2878] = 1'd0;
    assign memhint[2879] = 1'd0;
    assign memhint[2880] = 1'd0;
    assign memhint[2881] = 1'd0;
    assign memhint[2882] = 1'd0;
    assign memhint[2883] = 1'd0;
    assign memhint[2884] = 1'd0;
    assign memhint[2885] = 1'd0;
    assign memhint[2886] = 1'd0;
    assign memhint[2887] = 1'd0;
    assign memhint[2888] = 1'd0;
    assign memhint[2889] = 1'd0;
    assign memhint[2890] = 1'd0;
    assign memhint[2891] = 1'd0;
    assign memhint[2892] = 1'd0;
    assign memhint[2893] = 1'd0;
    assign memhint[2894] = 1'd0;
    assign memhint[2895] = 1'd0;
    assign memhint[2896] = 1'd1;
    assign memhint[2897] = 1'd1;
    assign memhint[2898] = 1'd0;
    assign memhint[2899] = 1'd0;
    assign memhint[2900] = 1'd0;
    assign memhint[2901] = 1'd0;
    assign memhint[2902] = 1'd0;
    assign memhint[2903] = 1'd0;
    assign memhint[2904] = 1'd0;
    assign memhint[2905] = 1'd0;
    assign memhint[2906] = 1'd0;
    assign memhint[2907] = 1'd0;
    assign memhint[2908] = 1'd0;
    assign memhint[2909] = 1'd0;
    assign memhint[2910] = 1'd0;
    assign memhint[2911] = 1'd0;
    assign memhint[2912] = 1'd0;
    assign memhint[2913] = 1'd1;
    assign memhint[2914] = 1'd1;
    assign memhint[2915] = 1'd0;
    assign memhint[2916] = 1'd0;
    assign memhint[2917] = 1'd0;
    assign memhint[2918] = 1'd0;
    assign memhint[2919] = 1'd0;
    assign memhint[2920] = 1'd0;
    assign memhint[2921] = 1'd0;
    assign memhint[2922] = 1'd0;
    assign memhint[2923] = 1'd0;
    assign memhint[2924] = 1'd0;
    assign memhint[2925] = 1'd1;
    assign memhint[2926] = 1'd1;
    assign memhint[2927] = 1'd0;
    assign memhint[2928] = 1'd0;
    assign memhint[2929] = 1'd0;
    assign memhint[2930] = 1'd0;
    assign memhint[2931] = 1'd0;
    assign memhint[2932] = 1'd1;
    assign memhint[2933] = 1'd1;
    assign memhint[2934] = 1'd0;
    assign memhint[2935] = 1'd0;
    assign memhint[2936] = 1'd0;
    assign memhint[2937] = 1'd0;
    assign memhint[2938] = 1'd0;
    assign memhint[2939] = 1'd0;
    assign memhint[2940] = 1'd0;
    assign memhint[2941] = 1'd0;
    assign memhint[2942] = 1'd0;
    assign memhint[2943] = 1'd0;
    assign memhint[2944] = 1'd0;
    assign memhint[2945] = 1'd0;
    assign memhint[2946] = 1'd0;
    assign memhint[2947] = 1'd0;
    assign memhint[2948] = 1'd0;
    assign memhint[2949] = 1'd0;
    assign memhint[2950] = 1'd0;
    assign memhint[2951] = 1'd0;
    assign memhint[2952] = 1'd1;
    assign memhint[2953] = 1'd1;
    assign memhint[2954] = 1'd0;
    assign memhint[2955] = 1'd0;
    assign memhint[2956] = 1'd0;
    assign memhint[2957] = 1'd1;
    assign memhint[2958] = 1'd1;
    assign memhint[2959] = 1'd0;
    assign memhint[2960] = 1'd0;
    assign memhint[2961] = 1'd0;
    assign memhint[2962] = 1'd0;
    assign memhint[2963] = 1'd0;
    assign memhint[2964] = 1'd0;
    assign memhint[2965] = 1'd0;
    assign memhint[2966] = 1'd0;
    assign memhint[2967] = 1'd0;
    assign memhint[2968] = 1'd0;
    assign memhint[2969] = 1'd0;
    assign memhint[2970] = 1'd0;
    assign memhint[2971] = 1'd0;
    assign memhint[2972] = 1'd1;
    assign memhint[2973] = 1'd1;
    assign memhint[2974] = 1'd1;
    assign memhint[2975] = 1'd0;
    assign memhint[2976] = 1'd0;
    assign memhint[2977] = 1'd1;
    assign memhint[2978] = 1'd1;
    assign memhint[2979] = 1'd1;
    assign memhint[2980] = 1'd0;
    assign memhint[2981] = 1'd0;
    assign memhint[2982] = 1'd0;
    assign memhint[2983] = 1'd0;
    assign memhint[2984] = 1'd0;
    assign memhint[2985] = 1'd0;
    assign memhint[2986] = 1'd1;
    assign memhint[2987] = 1'd1;
    assign memhint[2988] = 1'd1;
    assign memhint[2989] = 1'd0;
    assign memhint[2990] = 1'd0;
    assign memhint[2991] = 1'd0;
    assign memhint[2992] = 1'd0;
    assign memhint[2993] = 1'd0;
    assign memhint[2994] = 1'd0;
    assign memhint[2995] = 1'd0;
    assign memhint[2996] = 1'd0;
    assign memhint[2997] = 1'd0;
    assign memhint[2998] = 1'd0;
    assign memhint[2999] = 1'd0;
    assign memhint[3000] = 1'd0;
    assign memhint[3001] = 1'd0;
    assign memhint[3002] = 1'd1;
    assign memhint[3003] = 1'd1;
    assign memhint[3004] = 1'd0;
    assign memhint[3005] = 1'd0;
    assign memhint[3006] = 1'd0;
    assign memhint[3007] = 1'd0;
    assign memhint[3008] = 1'd0;
    assign memhint[3009] = 1'd0;
    assign memhint[3010] = 1'd0;
    assign memhint[3011] = 1'd0;
    assign memhint[3012] = 1'd0;
    assign memhint[3013] = 1'd0;
    assign memhint[3014] = 1'd0;
    assign memhint[3015] = 1'd0;
    assign memhint[3016] = 1'd0;
    assign memhint[3017] = 1'd0;
    assign memhint[3018] = 1'd0;
    assign memhint[3019] = 1'd1;
    assign memhint[3020] = 1'd1;
    assign memhint[3021] = 1'd0;
    assign memhint[3022] = 1'd0;
    assign memhint[3023] = 1'd0;
    assign memhint[3024] = 1'd0;
    assign memhint[3025] = 1'd0;
    assign memhint[3026] = 1'd0;
    assign memhint[3027] = 1'd0;
    assign memhint[3028] = 1'd0;
    assign memhint[3029] = 1'd0;
    assign memhint[3030] = 1'd0;
    assign memhint[3031] = 1'd0;
    assign memhint[3032] = 1'd0;
    assign memhint[3033] = 1'd0;
    assign memhint[3034] = 1'd1;
    assign memhint[3035] = 1'd1;
    assign memhint[3036] = 1'd0;
    assign memhint[3037] = 1'd0;
    assign memhint[3038] = 1'd0;
    assign memhint[3039] = 1'd0;
    assign memhint[3040] = 1'd0;
    assign memhint[3041] = 1'd0;
    assign memhint[3042] = 1'd0;
    assign memhint[3043] = 1'd0;
    assign memhint[3044] = 1'd0;
    assign memhint[3045] = 1'd0;
    assign memhint[3046] = 1'd0;
    assign memhint[3047] = 1'd0;
    assign memhint[3048] = 1'd0;
    assign memhint[3049] = 1'd0;
    assign memhint[3050] = 1'd1;
    assign memhint[3051] = 1'd1;
    assign memhint[3052] = 1'd0;
    assign memhint[3053] = 1'd0;
    assign memhint[3054] = 1'd0;
    assign memhint[3055] = 1'd0;
    assign memhint[3056] = 1'd0;
    assign memhint[3057] = 1'd0;
    assign memhint[3058] = 1'd0;
    assign memhint[3059] = 1'd0;
    assign memhint[3060] = 1'd0;
    assign memhint[3061] = 1'd0;
    assign memhint[3062] = 1'd0;
    assign memhint[3063] = 1'd0;
    assign memhint[3064] = 1'd0;
    assign memhint[3065] = 1'd0;
    assign memhint[3066] = 1'd0;
    assign memhint[3067] = 1'd0;
    assign memhint[3068] = 1'd0;
    assign memhint[3069] = 1'd0;
    assign memhint[3070] = 1'd0;
    assign memhint[3071] = 1'd0;
    assign memhint[3072] = 1'd0;
    assign memhint[3073] = 1'd0;
    assign memhint[3074] = 1'd0;
    assign memhint[3075] = 1'd0;
    assign memhint[3076] = 1'd0;
    assign memhint[3077] = 1'd0;
    assign memhint[3078] = 1'd0;
    assign memhint[3079] = 1'd1;
    assign memhint[3080] = 1'd1;
    assign memhint[3081] = 1'd0;
    assign memhint[3082] = 1'd0;
    assign memhint[3083] = 1'd0;
    assign memhint[3084] = 1'd0;
    assign memhint[3085] = 1'd0;
    assign memhint[3086] = 1'd0;
    assign memhint[3087] = 1'd0;
    assign memhint[3088] = 1'd0;
    assign memhint[3089] = 1'd0;
    assign memhint[3090] = 1'd0;
    assign memhint[3091] = 1'd0;
    assign memhint[3092] = 1'd0;
    assign memhint[3093] = 1'd0;
    assign memhint[3094] = 1'd0;
    assign memhint[3095] = 1'd0;
    assign memhint[3096] = 1'd0;
    assign memhint[3097] = 1'd0;
    assign memhint[3098] = 1'd0;
    assign memhint[3099] = 1'd0;
    assign memhint[3100] = 1'd0;
    assign memhint[3101] = 1'd0;
    assign memhint[3102] = 1'd0;
    assign memhint[3103] = 1'd1;
    assign memhint[3104] = 1'd1;
    assign memhint[3105] = 1'd0;
    assign memhint[3106] = 1'd0;
    assign memhint[3107] = 1'd0;
    assign memhint[3108] = 1'd0;
    assign memhint[3109] = 1'd0;
    assign memhint[3110] = 1'd1;
    assign memhint[3111] = 1'd1;
    assign memhint[3112] = 1'd0;
    assign memhint[3113] = 1'd0;
    assign memhint[3114] = 1'd0;
    assign memhint[3115] = 1'd0;
    assign memhint[3116] = 1'd0;
    assign memhint[3117] = 1'd0;
    assign memhint[3118] = 1'd0;
    assign memhint[3119] = 1'd0;
    assign memhint[3120] = 1'd0;
    assign memhint[3121] = 1'd0;
    assign memhint[3122] = 1'd0;
    assign memhint[3123] = 1'd0;
    assign memhint[3124] = 1'd0;
    assign memhint[3125] = 1'd0;
    assign memhint[3126] = 1'd0;
    assign memhint[3127] = 1'd0;
    assign memhint[3128] = 1'd0;
    assign memhint[3129] = 1'd0;
    assign memhint[3130] = 1'd0;
    assign memhint[3131] = 1'd1;
    assign memhint[3132] = 1'd1;
    assign memhint[3133] = 1'd1;
    assign memhint[3134] = 1'd0;
    assign memhint[3135] = 1'd0;
    assign memhint[3136] = 1'd0;
    assign memhint[3137] = 1'd0;
    assign memhint[3138] = 1'd0;
    assign memhint[3139] = 1'd0;
    assign memhint[3140] = 1'd0;
    assign memhint[3141] = 1'd0;
    assign memhint[3142] = 1'd0;
    assign memhint[3143] = 1'd0;
    assign memhint[3144] = 1'd0;
    assign memhint[3145] = 1'd0;
    assign memhint[3146] = 1'd1;
    assign memhint[3147] = 1'd1;
    assign memhint[3148] = 1'd0;
    assign memhint[3149] = 1'd0;
    assign memhint[3150] = 1'd0;
    assign memhint[3151] = 1'd0;
    assign memhint[3152] = 1'd0;
    assign memhint[3153] = 1'd0;
    assign memhint[3154] = 1'd0;
    assign memhint[3155] = 1'd0;
    assign memhint[3156] = 1'd0;
    assign memhint[3157] = 1'd0;
    assign memhint[3158] = 1'd0;
    assign memhint[3159] = 1'd0;
    assign memhint[3160] = 1'd0;
    assign memhint[3161] = 1'd0;
    assign memhint[3162] = 1'd0;
    assign memhint[3163] = 1'd0;
    assign memhint[3164] = 1'd0;
    assign memhint[3165] = 1'd0;
    assign memhint[3166] = 1'd0;
    assign memhint[3167] = 1'd0;
    assign memhint[3168] = 1'd1;
    assign memhint[3169] = 1'd1;
    assign memhint[3170] = 1'd0;
    assign memhint[3171] = 1'd0;
    assign memhint[3172] = 1'd0;
    assign memhint[3173] = 1'd0;
    assign memhint[3174] = 1'd0;
    assign memhint[3175] = 1'd1;
    assign memhint[3176] = 1'd1;
    assign memhint[3177] = 1'd0;
    assign memhint[3178] = 1'd0;
    assign memhint[3179] = 1'd0;
    assign memhint[3180] = 1'd1;
    assign memhint[3181] = 1'd1;
    assign memhint[3182] = 1'd1;
    assign memhint[3183] = 1'd0;
    assign memhint[3184] = 1'd0;
    assign memhint[3185] = 1'd0;
    assign memhint[3186] = 1'd0;
    assign memhint[3187] = 1'd0;
    assign memhint[3188] = 1'd0;
    assign memhint[3189] = 1'd0;
    assign memhint[3190] = 1'd0;
    assign memhint[3191] = 1'd1;
    assign memhint[3192] = 1'd1;
    assign memhint[3193] = 1'd0;
    assign memhint[3194] = 1'd0;
    assign memhint[3195] = 1'd0;
    assign memhint[3196] = 1'd0;
    assign memhint[3197] = 1'd0;
    assign memhint[3198] = 1'd1;
    assign memhint[3199] = 1'd1;
    assign memhint[3200] = 1'd1;
    assign memhint[3201] = 1'd0;
    assign memhint[3202] = 1'd0;
    assign memhint[3203] = 1'd0;
    assign memhint[3204] = 1'd0;
    assign memhint[3205] = 1'd0;
    assign memhint[3206] = 1'd0;
    assign memhint[3207] = 1'd0;
    assign memhint[3208] = 1'd0;
    assign memhint[3209] = 1'd0;
    assign memhint[3210] = 1'd0;
    assign memhint[3211] = 1'd0;
    assign memhint[3212] = 1'd0;
    assign memhint[3213] = 1'd0;
    assign memhint[3214] = 1'd0;
    assign memhint[3215] = 1'd0;
    assign memhint[3216] = 1'd0;
    assign memhint[3217] = 1'd0;
    assign memhint[3218] = 1'd0;
    assign memhint[3219] = 1'd0;
    assign memhint[3220] = 1'd0;
    assign memhint[3221] = 1'd0;
    assign memhint[3222] = 1'd0;
    assign memhint[3223] = 1'd0;
    assign memhint[3224] = 1'd0;
    assign memhint[3225] = 1'd0;
    assign memhint[3226] = 1'd0;
    assign memhint[3227] = 1'd0;
    assign memhint[3228] = 1'd0;
    assign memhint[3229] = 1'd0;
    assign memhint[3230] = 1'd0;
    assign memhint[3231] = 1'd0;
    assign memhint[3232] = 1'd0;
    assign memhint[3233] = 1'd0;
    assign memhint[3234] = 1'd0;
    assign memhint[3235] = 1'd0;
    assign memhint[3236] = 1'd0;
    assign memhint[3237] = 1'd0;
    assign memhint[3238] = 1'd1;
    assign memhint[3239] = 1'd1;
    assign memhint[3240] = 1'd0;
    assign memhint[3241] = 1'd0;
    assign memhint[3242] = 1'd0;
    assign memhint[3243] = 1'd0;
    assign memhint[3244] = 1'd0;
    assign memhint[3245] = 1'd0;
    assign memhint[3246] = 1'd0;
    assign memhint[3247] = 1'd0;
    assign memhint[3248] = 1'd1;
    assign memhint[3249] = 1'd1;
    assign memhint[3250] = 1'd0;
    assign memhint[3251] = 1'd0;
    assign memhint[3252] = 1'd0;
    assign memhint[3253] = 1'd0;
    assign memhint[3254] = 1'd0;
    assign memhint[3255] = 1'd0;
    assign memhint[3256] = 1'd0;
    assign memhint[3257] = 1'd0;
    assign memhint[3258] = 1'd0;
    assign memhint[3259] = 1'd0;
    assign memhint[3260] = 1'd0;
    assign memhint[3261] = 1'd0;
    assign memhint[3262] = 1'd0;
    assign memhint[3263] = 1'd0;
    assign memhint[3264] = 1'd0;
    assign memhint[3265] = 1'd0;
    assign memhint[3266] = 1'd0;
    assign memhint[3267] = 1'd0;
    assign memhint[3268] = 1'd0;
    assign memhint[3269] = 1'd0;
    assign memhint[3270] = 1'd1;
    assign memhint[3271] = 1'd1;
    assign memhint[3272] = 1'd0;
    assign memhint[3273] = 1'd0;
    assign memhint[3274] = 1'd0;
    assign memhint[3275] = 1'd0;
    assign memhint[3276] = 1'd0;
    assign memhint[3277] = 1'd0;
    assign memhint[3278] = 1'd0;
    assign memhint[3279] = 1'd0;
    assign memhint[3280] = 1'd0;
    assign memhint[3281] = 1'd0;
    assign memhint[3282] = 1'd0;
    assign memhint[3283] = 1'd0;
    assign memhint[3284] = 1'd0;
    assign memhint[3285] = 1'd0;
    assign memhint[3286] = 1'd1;
    assign memhint[3287] = 1'd1;
    assign memhint[3288] = 1'd0;
    assign memhint[3289] = 1'd0;
    assign memhint[3290] = 1'd0;
    assign memhint[3291] = 1'd0;
    assign memhint[3292] = 1'd0;
    assign memhint[3293] = 1'd0;
    assign memhint[3294] = 1'd0;
    assign memhint[3295] = 1'd0;
    assign memhint[3296] = 1'd0;
    assign memhint[3297] = 1'd1;
    assign memhint[3298] = 1'd1;
    assign memhint[3299] = 1'd1;
    assign memhint[3300] = 1'd0;
    assign memhint[3301] = 1'd0;
    assign memhint[3302] = 1'd0;
    assign memhint[3303] = 1'd0;
    assign memhint[3304] = 1'd0;
    assign memhint[3305] = 1'd1;
    assign memhint[3306] = 1'd1;
    assign memhint[3307] = 1'd0;
    assign memhint[3308] = 1'd0;
    assign memhint[3309] = 1'd0;
    assign memhint[3310] = 1'd0;
    assign memhint[3311] = 1'd0;
    assign memhint[3312] = 1'd0;
    assign memhint[3313] = 1'd0;
    assign memhint[3314] = 1'd0;
    assign memhint[3315] = 1'd0;
    assign memhint[3316] = 1'd0;
    assign memhint[3317] = 1'd0;
    assign memhint[3318] = 1'd0;
    assign memhint[3319] = 1'd0;
    assign memhint[3320] = 1'd0;
    assign memhint[3321] = 1'd0;
    assign memhint[3322] = 1'd0;
    assign memhint[3323] = 1'd0;
    assign memhint[3324] = 1'd1;
    assign memhint[3325] = 1'd1;
    assign memhint[3326] = 1'd0;
    assign memhint[3327] = 1'd0;
    assign memhint[3328] = 1'd0;
    assign memhint[3329] = 1'd0;
    assign memhint[3330] = 1'd0;
    assign memhint[3331] = 1'd1;
    assign memhint[3332] = 1'd1;
    assign memhint[3333] = 1'd0;
    assign memhint[3334] = 1'd0;
    assign memhint[3335] = 1'd0;
    assign memhint[3336] = 1'd0;
    assign memhint[3337] = 1'd0;
    assign memhint[3338] = 1'd0;
    assign memhint[3339] = 1'd0;
    assign memhint[3340] = 1'd0;
    assign memhint[3341] = 1'd0;
    assign memhint[3342] = 1'd0;
    assign memhint[3343] = 1'd0;
    assign memhint[3344] = 1'd0;
    assign memhint[3345] = 1'd0;
    assign memhint[3346] = 1'd1;
    assign memhint[3347] = 1'd1;
    assign memhint[3348] = 1'd0;
    assign memhint[3349] = 1'd0;
    assign memhint[3350] = 1'd1;
    assign memhint[3351] = 1'd1;
    assign memhint[3352] = 1'd0;
    assign memhint[3353] = 1'd0;
    assign memhint[3354] = 1'd0;
    assign memhint[3355] = 1'd0;
    assign memhint[3356] = 1'd0;
    assign memhint[3357] = 1'd0;
    assign memhint[3358] = 1'd0;
    assign memhint[3359] = 1'd0;
    assign memhint[3360] = 1'd1;
    assign memhint[3361] = 1'd1;
    assign memhint[3362] = 1'd1;
    assign memhint[3363] = 1'd1;
    assign memhint[3364] = 1'd0;
    assign memhint[3365] = 1'd0;
    assign memhint[3366] = 1'd0;
    assign memhint[3367] = 1'd0;
    assign memhint[3368] = 1'd0;
    assign memhint[3369] = 1'd0;
    assign memhint[3370] = 1'd0;
    assign memhint[3371] = 1'd0;
    assign memhint[3372] = 1'd0;
    assign memhint[3373] = 1'd0;
    assign memhint[3374] = 1'd0;
    assign memhint[3375] = 1'd1;
    assign memhint[3376] = 1'd1;
    assign memhint[3377] = 1'd1;
    assign memhint[3378] = 1'd1;
    assign memhint[3379] = 1'd1;
    assign memhint[3380] = 1'd1;
    assign memhint[3381] = 1'd1;
    assign memhint[3382] = 1'd1;
    assign memhint[3383] = 1'd1;
    assign memhint[3384] = 1'd1;
    assign memhint[3385] = 1'd1;
    assign memhint[3386] = 1'd1;
    assign memhint[3387] = 1'd1;
    assign memhint[3388] = 1'd0;
    assign memhint[3389] = 1'd0;
    assign memhint[3390] = 1'd0;
    assign memhint[3391] = 1'd0;
    assign memhint[3392] = 1'd1;
    assign memhint[3393] = 1'd1;
    assign memhint[3394] = 1'd0;
    assign memhint[3395] = 1'd0;
    assign memhint[3396] = 1'd0;
    assign memhint[3397] = 1'd0;
    assign memhint[3398] = 1'd0;
    assign memhint[3399] = 1'd0;
    assign memhint[3400] = 1'd0;
    assign memhint[3401] = 1'd0;
    assign memhint[3402] = 1'd0;
    assign memhint[3403] = 1'd0;
    assign memhint[3404] = 1'd0;
    assign memhint[3405] = 1'd0;
    assign memhint[3406] = 1'd0;
    assign memhint[3407] = 1'd1;
    assign memhint[3408] = 1'd1;
    assign memhint[3409] = 1'd1;
    assign memhint[3410] = 1'd1;
    assign memhint[3411] = 1'd1;
    assign memhint[3412] = 1'd1;
    assign memhint[3413] = 1'd1;
    assign memhint[3414] = 1'd1;
    assign memhint[3415] = 1'd1;
    assign memhint[3416] = 1'd1;
    assign memhint[3417] = 1'd1;
    assign memhint[3418] = 1'd1;
    assign memhint[3419] = 1'd1;
    assign memhint[3420] = 1'd0;
    assign memhint[3421] = 1'd0;
    assign memhint[3422] = 1'd0;
    assign memhint[3423] = 1'd1;
    assign memhint[3424] = 1'd1;
    assign memhint[3425] = 1'd0;
    assign memhint[3426] = 1'd0;
    assign memhint[3427] = 1'd0;
    assign memhint[3428] = 1'd0;
    assign memhint[3429] = 1'd0;
    assign memhint[3430] = 1'd0;
    assign memhint[3431] = 1'd0;
    assign memhint[3432] = 1'd0;
    assign memhint[3433] = 1'd0;
    assign memhint[3434] = 1'd0;
    assign memhint[3435] = 1'd0;
    assign memhint[3436] = 1'd0;
    assign memhint[3437] = 1'd0;
    assign memhint[3438] = 1'd0;
    assign memhint[3439] = 1'd0;
    assign memhint[3440] = 1'd0;
    assign memhint[3441] = 1'd0;
    assign memhint[3442] = 1'd0;
    assign memhint[3443] = 1'd0;
    assign memhint[3444] = 1'd0;
    assign memhint[3445] = 1'd0;
    assign memhint[3446] = 1'd0;
    assign memhint[3447] = 1'd0;
    assign memhint[3448] = 1'd0;
    assign memhint[3449] = 1'd0;
    assign memhint[3450] = 1'd0;
    assign memhint[3451] = 1'd0;
    assign memhint[3452] = 1'd1;
    assign memhint[3453] = 1'd1;
    assign memhint[3454] = 1'd0;
    assign memhint[3455] = 1'd0;
    assign memhint[3456] = 1'd0;
    assign memhint[3457] = 1'd0;
    assign memhint[3458] = 1'd0;
    assign memhint[3459] = 1'd0;
    assign memhint[3460] = 1'd0;
    assign memhint[3461] = 1'd0;
    assign memhint[3462] = 1'd0;
    assign memhint[3463] = 1'd0;
    assign memhint[3464] = 1'd0;
    assign memhint[3465] = 1'd0;
    assign memhint[3466] = 1'd0;
    assign memhint[3467] = 1'd0;
    assign memhint[3468] = 1'd0;
    assign memhint[3469] = 1'd0;
    assign memhint[3470] = 1'd0;
    assign memhint[3471] = 1'd0;
    assign memhint[3472] = 1'd0;
    assign memhint[3473] = 1'd0;
    assign memhint[3474] = 1'd0;
    assign memhint[3475] = 1'd0;
    assign memhint[3476] = 1'd1;
    assign memhint[3477] = 1'd1;
    assign memhint[3478] = 1'd0;
    assign memhint[3479] = 1'd0;
    assign memhint[3480] = 1'd0;
    assign memhint[3481] = 1'd0;
    assign memhint[3482] = 1'd0;
    assign memhint[3483] = 1'd1;
    assign memhint[3484] = 1'd1;
    assign memhint[3485] = 1'd0;
    assign memhint[3486] = 1'd0;
    assign memhint[3487] = 1'd0;
    assign memhint[3488] = 1'd0;
    assign memhint[3489] = 1'd0;
    assign memhint[3490] = 1'd0;
    assign memhint[3491] = 1'd0;
    assign memhint[3492] = 1'd0;
    assign memhint[3493] = 1'd0;
    assign memhint[3494] = 1'd0;
    assign memhint[3495] = 1'd0;
    assign memhint[3496] = 1'd0;
    assign memhint[3497] = 1'd0;
    assign memhint[3498] = 1'd0;
    assign memhint[3499] = 1'd0;
    assign memhint[3500] = 1'd0;
    assign memhint[3501] = 1'd0;
    assign memhint[3502] = 1'd0;
    assign memhint[3503] = 1'd0;
    assign memhint[3504] = 1'd0;
    assign memhint[3505] = 1'd1;
    assign memhint[3506] = 1'd1;
    assign memhint[3507] = 1'd1;
    assign memhint[3508] = 1'd1;
    assign memhint[3509] = 1'd0;
    assign memhint[3510] = 1'd0;
    assign memhint[3511] = 1'd0;
    assign memhint[3512] = 1'd0;
    assign memhint[3513] = 1'd0;
    assign memhint[3514] = 1'd0;
    assign memhint[3515] = 1'd0;
    assign memhint[3516] = 1'd0;
    assign memhint[3517] = 1'd0;
    assign memhint[3518] = 1'd0;
    assign memhint[3519] = 1'd1;
    assign memhint[3520] = 1'd1;
    assign memhint[3521] = 1'd0;
    assign memhint[3522] = 1'd0;
    assign memhint[3523] = 1'd0;
    assign memhint[3524] = 1'd0;
    assign memhint[3525] = 1'd0;
    assign memhint[3526] = 1'd0;
    assign memhint[3527] = 1'd0;
    assign memhint[3528] = 1'd0;
    assign memhint[3529] = 1'd0;
    assign memhint[3530] = 1'd0;
    assign memhint[3531] = 1'd0;
    assign memhint[3532] = 1'd0;
    assign memhint[3533] = 1'd0;
    assign memhint[3534] = 1'd0;
    assign memhint[3535] = 1'd0;
    assign memhint[3536] = 1'd0;
    assign memhint[3537] = 1'd0;
    assign memhint[3538] = 1'd0;
    assign memhint[3539] = 1'd0;
    assign memhint[3540] = 1'd0;
    assign memhint[3541] = 1'd1;
    assign memhint[3542] = 1'd1;
    assign memhint[3543] = 1'd0;
    assign memhint[3544] = 1'd0;
    assign memhint[3545] = 1'd0;
    assign memhint[3546] = 1'd0;
    assign memhint[3547] = 1'd0;
    assign memhint[3548] = 1'd1;
    assign memhint[3549] = 1'd1;
    assign memhint[3550] = 1'd0;
    assign memhint[3551] = 1'd0;
    assign memhint[3552] = 1'd0;
    assign memhint[3553] = 1'd0;
    assign memhint[3554] = 1'd1;
    assign memhint[3555] = 1'd1;
    assign memhint[3556] = 1'd0;
    assign memhint[3557] = 1'd0;
    assign memhint[3558] = 1'd0;
    assign memhint[3559] = 1'd0;
    assign memhint[3560] = 1'd0;
    assign memhint[3561] = 1'd0;
    assign memhint[3562] = 1'd0;
    assign memhint[3563] = 1'd0;
    assign memhint[3564] = 1'd1;
    assign memhint[3565] = 1'd1;
    assign memhint[3566] = 1'd0;
    assign memhint[3567] = 1'd0;
    assign memhint[3568] = 1'd0;
    assign memhint[3569] = 1'd0;
    assign memhint[3570] = 1'd0;
    assign memhint[3571] = 1'd1;
    assign memhint[3572] = 1'd1;
    assign memhint[3573] = 1'd0;
    assign memhint[3574] = 1'd0;
    assign memhint[3575] = 1'd0;
    assign memhint[3576] = 1'd0;
    assign memhint[3577] = 1'd0;
    assign memhint[3578] = 1'd0;
    assign memhint[3579] = 1'd0;
    assign memhint[3580] = 1'd0;
    assign memhint[3581] = 1'd0;
    assign memhint[3582] = 1'd0;
    assign memhint[3583] = 1'd0;
    assign memhint[3584] = 1'd0;
    assign memhint[3585] = 1'd0;
    assign memhint[3586] = 1'd0;
    assign memhint[3587] = 1'd0;
    assign memhint[3588] = 1'd0;
    assign memhint[3589] = 1'd0;
    assign memhint[3590] = 1'd0;
    assign memhint[3591] = 1'd0;
    assign memhint[3592] = 1'd0;
    assign memhint[3593] = 1'd0;
    assign memhint[3594] = 1'd0;
    assign memhint[3595] = 1'd0;
    assign memhint[3596] = 1'd0;
    assign memhint[3597] = 1'd0;
    assign memhint[3598] = 1'd0;
    assign memhint[3599] = 1'd0;
    assign memhint[3600] = 1'd0;
    assign memhint[3601] = 1'd0;
    assign memhint[3602] = 1'd0;
    assign memhint[3603] = 1'd0;
    assign memhint[3604] = 1'd0;
    assign memhint[3605] = 1'd0;
    assign memhint[3606] = 1'd0;
    assign memhint[3607] = 1'd0;
    assign memhint[3608] = 1'd0;
    assign memhint[3609] = 1'd0;
    assign memhint[3610] = 1'd0;
    assign memhint[3611] = 1'd1;
    assign memhint[3612] = 1'd1;
    assign memhint[3613] = 1'd0;
    assign memhint[3614] = 1'd0;
    assign memhint[3615] = 1'd0;
    assign memhint[3616] = 1'd0;
    assign memhint[3617] = 1'd0;
    assign memhint[3618] = 1'd0;
    assign memhint[3619] = 1'd0;
    assign memhint[3620] = 1'd0;
    assign memhint[3621] = 1'd1;
    assign memhint[3622] = 1'd1;
    assign memhint[3623] = 1'd0;
    assign memhint[3624] = 1'd0;
    assign memhint[3625] = 1'd0;
    assign memhint[3626] = 1'd0;
    assign memhint[3627] = 1'd0;
    assign memhint[3628] = 1'd0;
    assign memhint[3629] = 1'd0;
    assign memhint[3630] = 1'd0;
    assign memhint[3631] = 1'd0;
    assign memhint[3632] = 1'd0;
    assign memhint[3633] = 1'd0;
    assign memhint[3634] = 1'd0;
    assign memhint[3635] = 1'd0;
    assign memhint[3636] = 1'd0;
    assign memhint[3637] = 1'd0;
    assign memhint[3638] = 1'd0;
    assign memhint[3639] = 1'd0;
    assign memhint[3640] = 1'd0;
    assign memhint[3641] = 1'd0;
    assign memhint[3642] = 1'd0;
    assign memhint[3643] = 1'd1;
    assign memhint[3644] = 1'd1;
    assign memhint[3645] = 1'd0;
    assign memhint[3646] = 1'd0;
    assign memhint[3647] = 1'd0;
    assign memhint[3648] = 1'd0;
    assign memhint[3649] = 1'd0;
    assign memhint[3650] = 1'd0;
    assign memhint[3651] = 1'd0;
    assign memhint[3652] = 1'd0;
    assign memhint[3653] = 1'd0;
    assign memhint[3654] = 1'd0;
    assign memhint[3655] = 1'd0;
    assign memhint[3656] = 1'd0;
    assign memhint[3657] = 1'd0;
    assign memhint[3658] = 1'd0;
    assign memhint[3659] = 1'd1;
    assign memhint[3660] = 1'd1;
    assign memhint[3661] = 1'd0;
    assign memhint[3662] = 1'd0;
    assign memhint[3663] = 1'd0;
    assign memhint[3664] = 1'd0;
    assign memhint[3665] = 1'd0;
    assign memhint[3666] = 1'd0;
    assign memhint[3667] = 1'd0;
    assign memhint[3668] = 1'd0;
    assign memhint[3669] = 1'd1;
    assign memhint[3670] = 1'd1;
    assign memhint[3671] = 1'd1;
    assign memhint[3672] = 1'd0;
    assign memhint[3673] = 1'd0;
    assign memhint[3674] = 1'd0;
    assign memhint[3675] = 1'd0;
    assign memhint[3676] = 1'd0;
    assign memhint[3677] = 1'd0;
    assign memhint[3678] = 1'd1;
    assign memhint[3679] = 1'd1;
    assign memhint[3680] = 1'd0;
    assign memhint[3681] = 1'd0;
    assign memhint[3682] = 1'd0;
    assign memhint[3683] = 1'd0;
    assign memhint[3684] = 1'd0;
    assign memhint[3685] = 1'd0;
    assign memhint[3686] = 1'd0;
    assign memhint[3687] = 1'd0;
    assign memhint[3688] = 1'd0;
    assign memhint[3689] = 1'd0;
    assign memhint[3690] = 1'd0;
    assign memhint[3691] = 1'd0;
    assign memhint[3692] = 1'd0;
    assign memhint[3693] = 1'd0;
    assign memhint[3694] = 1'd0;
    assign memhint[3695] = 1'd0;
    assign memhint[3696] = 1'd0;
    assign memhint[3697] = 1'd1;
    assign memhint[3698] = 1'd1;
    assign memhint[3699] = 1'd0;
    assign memhint[3700] = 1'd0;
    assign memhint[3701] = 1'd0;
    assign memhint[3702] = 1'd0;
    assign memhint[3703] = 1'd0;
    assign memhint[3704] = 1'd1;
    assign memhint[3705] = 1'd1;
    assign memhint[3706] = 1'd0;
    assign memhint[3707] = 1'd0;
    assign memhint[3708] = 1'd0;
    assign memhint[3709] = 1'd0;
    assign memhint[3710] = 1'd0;
    assign memhint[3711] = 1'd0;
    assign memhint[3712] = 1'd0;
    assign memhint[3713] = 1'd0;
    assign memhint[3714] = 1'd0;
    assign memhint[3715] = 1'd0;
    assign memhint[3716] = 1'd0;
    assign memhint[3717] = 1'd0;
    assign memhint[3718] = 1'd0;
    assign memhint[3719] = 1'd0;
    assign memhint[3720] = 1'd1;
    assign memhint[3721] = 1'd1;
    assign memhint[3722] = 1'd1;
    assign memhint[3723] = 1'd1;
    assign memhint[3724] = 1'd0;
    assign memhint[3725] = 1'd0;
    assign memhint[3726] = 1'd0;
    assign memhint[3727] = 1'd0;
    assign memhint[3728] = 1'd0;
    assign memhint[3729] = 1'd0;
    assign memhint[3730] = 1'd0;
    assign memhint[3731] = 1'd0;
    assign memhint[3732] = 1'd0;
    assign memhint[3733] = 1'd0;
    assign memhint[3734] = 1'd0;
    assign memhint[3735] = 1'd1;
    assign memhint[3736] = 1'd1;
    assign memhint[3737] = 1'd1;
    assign memhint[3738] = 1'd0;
    assign memhint[3739] = 1'd0;
    assign memhint[3740] = 1'd0;
    assign memhint[3741] = 1'd0;
    assign memhint[3742] = 1'd0;
    assign memhint[3743] = 1'd0;
    assign memhint[3744] = 1'd0;
    assign memhint[3745] = 1'd0;
    assign memhint[3746] = 1'd0;
    assign memhint[3747] = 1'd0;
    assign memhint[3748] = 1'd1;
    assign memhint[3749] = 1'd1;
    assign memhint[3750] = 1'd1;
    assign memhint[3751] = 1'd1;
    assign memhint[3752] = 1'd1;
    assign memhint[3753] = 1'd1;
    assign memhint[3754] = 1'd1;
    assign memhint[3755] = 1'd1;
    assign memhint[3756] = 1'd1;
    assign memhint[3757] = 1'd1;
    assign memhint[3758] = 1'd1;
    assign memhint[3759] = 1'd1;
    assign memhint[3760] = 1'd1;
    assign memhint[3761] = 1'd0;
    assign memhint[3762] = 1'd0;
    assign memhint[3763] = 1'd0;
    assign memhint[3764] = 1'd0;
    assign memhint[3765] = 1'd1;
    assign memhint[3766] = 1'd1;
    assign memhint[3767] = 1'd0;
    assign memhint[3768] = 1'd0;
    assign memhint[3769] = 1'd0;
    assign memhint[3770] = 1'd0;
    assign memhint[3771] = 1'd0;
    assign memhint[3772] = 1'd0;
    assign memhint[3773] = 1'd0;
    assign memhint[3774] = 1'd0;
    assign memhint[3775] = 1'd0;
    assign memhint[3776] = 1'd0;
    assign memhint[3777] = 1'd0;
    assign memhint[3778] = 1'd0;
    assign memhint[3779] = 1'd0;
    assign memhint[3780] = 1'd1;
    assign memhint[3781] = 1'd1;
    assign memhint[3782] = 1'd1;
    assign memhint[3783] = 1'd1;
    assign memhint[3784] = 1'd1;
    assign memhint[3785] = 1'd1;
    assign memhint[3786] = 1'd1;
    assign memhint[3787] = 1'd1;
    assign memhint[3788] = 1'd1;
    assign memhint[3789] = 1'd1;
    assign memhint[3790] = 1'd1;
    assign memhint[3791] = 1'd1;
    assign memhint[3792] = 1'd1;
    assign memhint[3793] = 1'd0;
    assign memhint[3794] = 1'd0;
    assign memhint[3795] = 1'd0;
    assign memhint[3796] = 1'd1;
    assign memhint[3797] = 1'd1;
    assign memhint[3798] = 1'd0;
    assign memhint[3799] = 1'd0;
    assign memhint[3800] = 1'd0;
    assign memhint[3801] = 1'd0;
    assign memhint[3802] = 1'd0;
    assign memhint[3803] = 1'd0;
    assign memhint[3804] = 1'd0;
    assign memhint[3805] = 1'd0;
    assign memhint[3806] = 1'd0;
    assign memhint[3807] = 1'd0;
    assign memhint[3808] = 1'd0;
    assign memhint[3809] = 1'd0;
    assign memhint[3810] = 1'd0;
    assign memhint[3811] = 1'd0;
    assign memhint[3812] = 1'd0;
    assign memhint[3813] = 1'd0;
    assign memhint[3814] = 1'd0;
    assign memhint[3815] = 1'd0;
    assign memhint[3816] = 1'd0;
    assign memhint[3817] = 1'd0;
    assign memhint[3818] = 1'd0;
    assign memhint[3819] = 1'd0;
    assign memhint[3820] = 1'd0;
    assign memhint[3821] = 1'd0;
    assign memhint[3822] = 1'd0;
    assign memhint[3823] = 1'd0;
    assign memhint[3824] = 1'd0;
    assign memhint[3825] = 1'd1;
    assign memhint[3826] = 1'd1;
    assign memhint[3827] = 1'd0;
    assign memhint[3828] = 1'd0;
    assign memhint[3829] = 1'd0;
    assign memhint[3830] = 1'd0;
    assign memhint[3831] = 1'd0;
    assign memhint[3832] = 1'd0;
    assign memhint[3833] = 1'd0;
    assign memhint[3834] = 1'd0;
    assign memhint[3835] = 1'd0;
    assign memhint[3836] = 1'd0;
    assign memhint[3837] = 1'd0;
    assign memhint[3838] = 1'd0;
    assign memhint[3839] = 1'd0;
    assign memhint[3840] = 1'd0;
    assign memhint[3841] = 1'd0;
    assign memhint[3842] = 1'd0;
    assign memhint[3843] = 1'd0;
    assign memhint[3844] = 1'd0;
    assign memhint[3845] = 1'd0;
    assign memhint[3846] = 1'd0;
    assign memhint[3847] = 1'd0;
    assign memhint[3848] = 1'd1;
    assign memhint[3849] = 1'd1;
    assign memhint[3850] = 1'd1;
    assign memhint[3851] = 1'd0;
    assign memhint[3852] = 1'd0;
    assign memhint[3853] = 1'd0;
    assign memhint[3854] = 1'd0;
    assign memhint[3855] = 1'd0;
    assign memhint[3856] = 1'd1;
    assign memhint[3857] = 1'd1;
    assign memhint[3858] = 1'd1;
    assign memhint[3859] = 1'd0;
    assign memhint[3860] = 1'd0;
    assign memhint[3861] = 1'd0;
    assign memhint[3862] = 1'd0;
    assign memhint[3863] = 1'd0;
    assign memhint[3864] = 1'd0;
    assign memhint[3865] = 1'd0;
    assign memhint[3866] = 1'd0;
    assign memhint[3867] = 1'd0;
    assign memhint[3868] = 1'd0;
    assign memhint[3869] = 1'd0;
    assign memhint[3870] = 1'd0;
    assign memhint[3871] = 1'd0;
    assign memhint[3872] = 1'd0;
    assign memhint[3873] = 1'd0;
    assign memhint[3874] = 1'd0;
    assign memhint[3875] = 1'd0;
    assign memhint[3876] = 1'd0;
    assign memhint[3877] = 1'd0;
    assign memhint[3878] = 1'd0;
    assign memhint[3879] = 1'd0;
    assign memhint[3880] = 1'd1;
    assign memhint[3881] = 1'd1;
    assign memhint[3882] = 1'd1;
    assign memhint[3883] = 1'd0;
    assign memhint[3884] = 1'd0;
    assign memhint[3885] = 1'd0;
    assign memhint[3886] = 1'd0;
    assign memhint[3887] = 1'd0;
    assign memhint[3888] = 1'd0;
    assign memhint[3889] = 1'd0;
    assign memhint[3890] = 1'd0;
    assign memhint[3891] = 1'd0;
    assign memhint[3892] = 1'd1;
    assign memhint[3893] = 1'd1;
    assign memhint[3894] = 1'd0;
    assign memhint[3895] = 1'd0;
    assign memhint[3896] = 1'd0;
    assign memhint[3897] = 1'd0;
    assign memhint[3898] = 1'd0;
    assign memhint[3899] = 1'd0;
    assign memhint[3900] = 1'd0;
    assign memhint[3901] = 1'd0;
    assign memhint[3902] = 1'd0;
    assign memhint[3903] = 1'd0;
    assign memhint[3904] = 1'd0;
    assign memhint[3905] = 1'd0;
    assign memhint[3906] = 1'd0;
    assign memhint[3907] = 1'd0;
    assign memhint[3908] = 1'd0;
    assign memhint[3909] = 1'd0;
    assign memhint[3910] = 1'd0;
    assign memhint[3911] = 1'd0;
    assign memhint[3912] = 1'd0;
    assign memhint[3913] = 1'd0;
    assign memhint[3914] = 1'd1;
    assign memhint[3915] = 1'd1;
    assign memhint[3916] = 1'd0;
    assign memhint[3917] = 1'd0;
    assign memhint[3918] = 1'd0;
    assign memhint[3919] = 1'd0;
    assign memhint[3920] = 1'd0;
    assign memhint[3921] = 1'd1;
    assign memhint[3922] = 1'd1;
    assign memhint[3923] = 1'd0;
    assign memhint[3924] = 1'd0;
    assign memhint[3925] = 1'd0;
    assign memhint[3926] = 1'd0;
    assign memhint[3927] = 1'd0;
    assign memhint[3928] = 1'd1;
    assign memhint[3929] = 1'd1;
    assign memhint[3930] = 1'd0;
    assign memhint[3931] = 1'd0;
    assign memhint[3932] = 1'd0;
    assign memhint[3933] = 1'd0;
    assign memhint[3934] = 1'd0;
    assign memhint[3935] = 1'd0;
    assign memhint[3936] = 1'd0;
    assign memhint[3937] = 1'd1;
    assign memhint[3938] = 1'd1;
    assign memhint[3939] = 1'd0;
    assign memhint[3940] = 1'd0;
    assign memhint[3941] = 1'd0;
    assign memhint[3942] = 1'd0;
    assign memhint[3943] = 1'd0;
    assign memhint[3944] = 1'd1;
    assign memhint[3945] = 1'd1;
    assign memhint[3946] = 1'd0;
    assign memhint[3947] = 1'd0;
    assign memhint[3948] = 1'd0;
    assign memhint[3949] = 1'd0;
    assign memhint[3950] = 1'd0;
    assign memhint[3951] = 1'd0;
    assign memhint[3952] = 1'd0;
    assign memhint[3953] = 1'd0;
    assign memhint[3954] = 1'd0;
    assign memhint[3955] = 1'd0;
    assign memhint[3956] = 1'd0;
    assign memhint[3957] = 1'd0;
    assign memhint[3958] = 1'd0;
    assign memhint[3959] = 1'd0;
    assign memhint[3960] = 1'd0;
    assign memhint[3961] = 1'd0;
    assign memhint[3962] = 1'd0;
    assign memhint[3963] = 1'd0;
    assign memhint[3964] = 1'd0;
    assign memhint[3965] = 1'd0;
    assign memhint[3966] = 1'd0;
    assign memhint[3967] = 1'd0;
    assign memhint[3968] = 1'd0;
    assign memhint[3969] = 1'd0;
    assign memhint[3970] = 1'd0;
    assign memhint[3971] = 1'd0;
    assign memhint[3972] = 1'd0;
    assign memhint[3973] = 1'd0;
    assign memhint[3974] = 1'd0;
    assign memhint[3975] = 1'd0;
    assign memhint[3976] = 1'd0;
    assign memhint[3977] = 1'd0;
    assign memhint[3978] = 1'd0;
    assign memhint[3979] = 1'd0;
    assign memhint[3980] = 1'd0;
    assign memhint[3981] = 1'd0;
    assign memhint[3982] = 1'd0;
    assign memhint[3983] = 1'd0;
    assign memhint[3984] = 1'd1;
    assign memhint[3985] = 1'd1;
    assign memhint[3986] = 1'd0;
    assign memhint[3987] = 1'd0;
    assign memhint[3988] = 1'd0;
    assign memhint[3989] = 1'd0;
    assign memhint[3990] = 1'd0;
    assign memhint[3991] = 1'd0;
    assign memhint[3992] = 1'd0;
    assign memhint[3993] = 1'd0;
    assign memhint[3994] = 1'd1;
    assign memhint[3995] = 1'd1;
    assign memhint[3996] = 1'd0;
    assign memhint[3997] = 1'd0;
    assign memhint[3998] = 1'd0;
    assign memhint[3999] = 1'd0;
    assign memhint[4000] = 1'd0;
    assign memhint[4001] = 1'd0;
    assign memhint[4002] = 1'd0;
    assign memhint[4003] = 1'd0;
    assign memhint[4004] = 1'd0;
    assign memhint[4005] = 1'd0;
    assign memhint[4006] = 1'd0;
    assign memhint[4007] = 1'd0;
    assign memhint[4008] = 1'd0;
    assign memhint[4009] = 1'd0;
    assign memhint[4010] = 1'd0;
    assign memhint[4011] = 1'd0;
    assign memhint[4012] = 1'd0;
    assign memhint[4013] = 1'd0;
    assign memhint[4014] = 1'd0;
    assign memhint[4015] = 1'd0;
    assign memhint[4016] = 1'd1;
    assign memhint[4017] = 1'd1;
    assign memhint[4018] = 1'd0;
    assign memhint[4019] = 1'd0;
    assign memhint[4020] = 1'd0;
    assign memhint[4021] = 1'd0;
    assign memhint[4022] = 1'd0;
    assign memhint[4023] = 1'd0;
    assign memhint[4024] = 1'd0;
    assign memhint[4025] = 1'd0;
    assign memhint[4026] = 1'd0;
    assign memhint[4027] = 1'd0;
    assign memhint[4028] = 1'd0;
    assign memhint[4029] = 1'd0;
    assign memhint[4030] = 1'd0;
    assign memhint[4031] = 1'd0;
    assign memhint[4032] = 1'd1;
    assign memhint[4033] = 1'd1;
    assign memhint[4034] = 1'd1;
    assign memhint[4035] = 1'd1;
    assign memhint[4036] = 1'd1;
    assign memhint[4037] = 1'd1;
    assign memhint[4038] = 1'd1;
    assign memhint[4039] = 1'd1;
    assign memhint[4040] = 1'd1;
    assign memhint[4041] = 1'd1;
    assign memhint[4042] = 1'd1;
    assign memhint[4043] = 1'd1;
    assign memhint[4044] = 1'd0;
    assign memhint[4045] = 1'd0;
    assign memhint[4046] = 1'd0;
    assign memhint[4047] = 1'd0;
    assign memhint[4048] = 1'd0;
    assign memhint[4049] = 1'd0;
    assign memhint[4050] = 1'd0;
    assign memhint[4051] = 1'd1;
    assign memhint[4052] = 1'd1;
    assign memhint[4053] = 1'd0;
    assign memhint[4054] = 1'd0;
    assign memhint[4055] = 1'd0;
    assign memhint[4056] = 1'd0;
    assign memhint[4057] = 1'd0;
    assign memhint[4058] = 1'd0;
    assign memhint[4059] = 1'd0;
    assign memhint[4060] = 1'd0;
    assign memhint[4061] = 1'd0;
    assign memhint[4062] = 1'd0;
    assign memhint[4063] = 1'd0;
    assign memhint[4064] = 1'd0;
    assign memhint[4065] = 1'd0;
    assign memhint[4066] = 1'd0;
    assign memhint[4067] = 1'd0;
    assign memhint[4068] = 1'd0;
    assign memhint[4069] = 1'd1;
    assign memhint[4070] = 1'd1;
    assign memhint[4071] = 1'd1;
    assign memhint[4072] = 1'd0;
    assign memhint[4073] = 1'd0;
    assign memhint[4074] = 1'd0;
    assign memhint[4075] = 1'd0;
    assign memhint[4076] = 1'd0;
    assign memhint[4077] = 1'd1;
    assign memhint[4078] = 1'd1;
    assign memhint[4079] = 1'd1;
    assign memhint[4080] = 1'd0;
    assign memhint[4081] = 1'd0;
    assign memhint[4082] = 1'd0;
    assign memhint[4083] = 1'd0;
    assign memhint[4084] = 1'd0;
    assign memhint[4085] = 1'd0;
    assign memhint[4086] = 1'd0;
    assign memhint[4087] = 1'd0;
    assign memhint[4088] = 1'd0;
    assign memhint[4089] = 1'd0;
    assign memhint[4090] = 1'd0;
    assign memhint[4091] = 1'd0;
    assign memhint[4092] = 1'd0;
    assign memhint[4093] = 1'd1;
    assign memhint[4094] = 1'd1;
    assign memhint[4095] = 1'd1;
    assign memhint[4096] = 1'd1;
    assign memhint[4097] = 1'd0;
    assign memhint[4098] = 1'd0;
    assign memhint[4099] = 1'd0;
    assign memhint[4100] = 1'd0;
    assign memhint[4101] = 1'd0;
    assign memhint[4102] = 1'd0;
    assign memhint[4103] = 1'd0;
    assign memhint[4104] = 1'd0;
    assign memhint[4105] = 1'd0;
    assign memhint[4106] = 1'd0;
    assign memhint[4107] = 1'd0;
    assign memhint[4108] = 1'd0;
    assign memhint[4109] = 1'd1;
    assign memhint[4110] = 1'd1;
    assign memhint[4111] = 1'd1;
    assign memhint[4112] = 1'd1;
    assign memhint[4113] = 1'd0;
    assign memhint[4114] = 1'd0;
    assign memhint[4115] = 1'd0;
    assign memhint[4116] = 1'd0;
    assign memhint[4117] = 1'd0;
    assign memhint[4118] = 1'd0;
    assign memhint[4119] = 1'd0;
    assign memhint[4120] = 1'd0;
    assign memhint[4121] = 1'd1;
    assign memhint[4122] = 1'd1;
    assign memhint[4123] = 1'd0;
    assign memhint[4124] = 1'd0;
    assign memhint[4125] = 1'd0;
    assign memhint[4126] = 1'd0;
    assign memhint[4127] = 1'd0;
    assign memhint[4128] = 1'd0;
    assign memhint[4129] = 1'd0;
    assign memhint[4130] = 1'd0;
    assign memhint[4131] = 1'd0;
    assign memhint[4132] = 1'd0;
    assign memhint[4133] = 1'd0;
    assign memhint[4134] = 1'd0;
    assign memhint[4135] = 1'd0;
    assign memhint[4136] = 1'd0;
    assign memhint[4137] = 1'd0;
    assign memhint[4138] = 1'd1;
    assign memhint[4139] = 1'd1;
    assign memhint[4140] = 1'd0;
    assign memhint[4141] = 1'd0;
    assign memhint[4142] = 1'd0;
    assign memhint[4143] = 1'd0;
    assign memhint[4144] = 1'd0;
    assign memhint[4145] = 1'd0;
    assign memhint[4146] = 1'd0;
    assign memhint[4147] = 1'd0;
    assign memhint[4148] = 1'd0;
    assign memhint[4149] = 1'd0;
    assign memhint[4150] = 1'd0;
    assign memhint[4151] = 1'd0;
    assign memhint[4152] = 1'd0;
    assign memhint[4153] = 1'd1;
    assign memhint[4154] = 1'd1;
    assign memhint[4155] = 1'd0;
    assign memhint[4156] = 1'd0;
    assign memhint[4157] = 1'd0;
    assign memhint[4158] = 1'd0;
    assign memhint[4159] = 1'd0;
    assign memhint[4160] = 1'd0;
    assign memhint[4161] = 1'd0;
    assign memhint[4162] = 1'd0;
    assign memhint[4163] = 1'd0;
    assign memhint[4164] = 1'd0;
    assign memhint[4165] = 1'd0;
    assign memhint[4166] = 1'd0;
    assign memhint[4167] = 1'd0;
    assign memhint[4168] = 1'd0;
    assign memhint[4169] = 1'd1;
    assign memhint[4170] = 1'd1;
    assign memhint[4171] = 1'd0;
    assign memhint[4172] = 1'd0;
    assign memhint[4173] = 1'd0;
    assign memhint[4174] = 1'd0;
    assign memhint[4175] = 1'd0;
    assign memhint[4176] = 1'd0;
    assign memhint[4177] = 1'd0;
    assign memhint[4178] = 1'd0;
    assign memhint[4179] = 1'd0;
    assign memhint[4180] = 1'd0;
    assign memhint[4181] = 1'd0;
    assign memhint[4182] = 1'd0;
    assign memhint[4183] = 1'd0;
    assign memhint[4184] = 1'd0;
    assign memhint[4185] = 1'd0;
    assign memhint[4186] = 1'd0;
    assign memhint[4187] = 1'd0;
    assign memhint[4188] = 1'd0;
    assign memhint[4189] = 1'd0;
    assign memhint[4190] = 1'd0;
    assign memhint[4191] = 1'd0;
    assign memhint[4192] = 1'd0;
    assign memhint[4193] = 1'd0;
    assign memhint[4194] = 1'd0;
    assign memhint[4195] = 1'd0;
    assign memhint[4196] = 1'd0;
    assign memhint[4197] = 1'd0;
    assign memhint[4198] = 1'd1;
    assign memhint[4199] = 1'd1;
    assign memhint[4200] = 1'd0;
    assign memhint[4201] = 1'd0;
    assign memhint[4202] = 1'd0;
    assign memhint[4203] = 1'd0;
    assign memhint[4204] = 1'd0;
    assign memhint[4205] = 1'd0;
    assign memhint[4206] = 1'd0;
    assign memhint[4207] = 1'd0;
    assign memhint[4208] = 1'd0;
    assign memhint[4209] = 1'd0;
    assign memhint[4210] = 1'd0;
    assign memhint[4211] = 1'd0;
    assign memhint[4212] = 1'd0;
    assign memhint[4213] = 1'd0;
    assign memhint[4214] = 1'd0;
    assign memhint[4215] = 1'd0;
    assign memhint[4216] = 1'd0;
    assign memhint[4217] = 1'd0;
    assign memhint[4218] = 1'd0;
    assign memhint[4219] = 1'd0;
    assign memhint[4220] = 1'd0;
    assign memhint[4221] = 1'd1;
    assign memhint[4222] = 1'd1;
    assign memhint[4223] = 1'd0;
    assign memhint[4224] = 1'd0;
    assign memhint[4225] = 1'd0;
    assign memhint[4226] = 1'd0;
    assign memhint[4227] = 1'd0;
    assign memhint[4228] = 1'd0;
    assign memhint[4229] = 1'd0;
    assign memhint[4230] = 1'd1;
    assign memhint[4231] = 1'd1;
    assign memhint[4232] = 1'd0;
    assign memhint[4233] = 1'd0;
    assign memhint[4234] = 1'd0;
    assign memhint[4235] = 1'd0;
    assign memhint[4236] = 1'd0;
    assign memhint[4237] = 1'd0;
    assign memhint[4238] = 1'd0;
    assign memhint[4239] = 1'd0;
    assign memhint[4240] = 1'd0;
    assign memhint[4241] = 1'd0;
    assign memhint[4242] = 1'd0;
    assign memhint[4243] = 1'd0;
    assign memhint[4244] = 1'd0;
    assign memhint[4245] = 1'd0;
    assign memhint[4246] = 1'd0;
    assign memhint[4247] = 1'd0;
    assign memhint[4248] = 1'd0;
    assign memhint[4249] = 1'd0;
    assign memhint[4250] = 1'd0;
    assign memhint[4251] = 1'd0;
    assign memhint[4252] = 1'd0;
    assign memhint[4253] = 1'd0;
    assign memhint[4254] = 1'd1;
    assign memhint[4255] = 1'd1;
    assign memhint[4256] = 1'd1;
    assign memhint[4257] = 1'd1;
    assign memhint[4258] = 1'd0;
    assign memhint[4259] = 1'd0;
    assign memhint[4260] = 1'd0;
    assign memhint[4261] = 1'd0;
    assign memhint[4262] = 1'd0;
    assign memhint[4263] = 1'd0;
    assign memhint[4264] = 1'd0;
    assign memhint[4265] = 1'd1;
    assign memhint[4266] = 1'd1;
    assign memhint[4267] = 1'd0;
    assign memhint[4268] = 1'd0;
    assign memhint[4269] = 1'd0;
    assign memhint[4270] = 1'd0;
    assign memhint[4271] = 1'd0;
    assign memhint[4272] = 1'd0;
    assign memhint[4273] = 1'd0;
    assign memhint[4274] = 1'd0;
    assign memhint[4275] = 1'd0;
    assign memhint[4276] = 1'd0;
    assign memhint[4277] = 1'd0;
    assign memhint[4278] = 1'd0;
    assign memhint[4279] = 1'd0;
    assign memhint[4280] = 1'd0;
    assign memhint[4281] = 1'd0;
    assign memhint[4282] = 1'd0;
    assign memhint[4283] = 1'd0;
    assign memhint[4284] = 1'd0;
    assign memhint[4285] = 1'd0;
    assign memhint[4286] = 1'd0;
    assign memhint[4287] = 1'd1;
    assign memhint[4288] = 1'd1;
    assign memhint[4289] = 1'd0;
    assign memhint[4290] = 1'd0;
    assign memhint[4291] = 1'd0;
    assign memhint[4292] = 1'd0;
    assign memhint[4293] = 1'd0;
    assign memhint[4294] = 1'd1;
    assign memhint[4295] = 1'd1;
    assign memhint[4296] = 1'd0;
    assign memhint[4297] = 1'd0;
    assign memhint[4298] = 1'd0;
    assign memhint[4299] = 1'd0;
    assign memhint[4300] = 1'd0;
    assign memhint[4301] = 1'd0;
    assign memhint[4302] = 1'd1;
    assign memhint[4303] = 1'd1;
    assign memhint[4304] = 1'd0;
    assign memhint[4305] = 1'd0;
    assign memhint[4306] = 1'd0;
    assign memhint[4307] = 1'd0;
    assign memhint[4308] = 1'd0;
    assign memhint[4309] = 1'd0;
    assign memhint[4310] = 1'd1;
    assign memhint[4311] = 1'd1;
    assign memhint[4312] = 1'd0;
    assign memhint[4313] = 1'd0;
    assign memhint[4314] = 1'd0;
    assign memhint[4315] = 1'd0;
    assign memhint[4316] = 1'd0;
    assign memhint[4317] = 1'd1;
    assign memhint[4318] = 1'd1;
    assign memhint[4319] = 1'd0;
    assign memhint[4320] = 1'd0;
    assign memhint[4321] = 1'd0;
    assign memhint[4322] = 1'd0;
    assign memhint[4323] = 1'd0;
    assign memhint[4324] = 1'd0;
    assign memhint[4325] = 1'd0;
    assign memhint[4326] = 1'd0;
    assign memhint[4327] = 1'd0;
    assign memhint[4328] = 1'd0;
    assign memhint[4329] = 1'd0;
    assign memhint[4330] = 1'd0;
    assign memhint[4331] = 1'd0;
    assign memhint[4332] = 1'd0;
    assign memhint[4333] = 1'd0;
    assign memhint[4334] = 1'd0;
    assign memhint[4335] = 1'd0;
    assign memhint[4336] = 1'd0;
    assign memhint[4337] = 1'd0;
    assign memhint[4338] = 1'd0;
    assign memhint[4339] = 1'd0;
    assign memhint[4340] = 1'd0;
    assign memhint[4341] = 1'd0;
    assign memhint[4342] = 1'd0;
    assign memhint[4343] = 1'd0;
    assign memhint[4344] = 1'd0;
    assign memhint[4345] = 1'd0;
    assign memhint[4346] = 1'd0;
    assign memhint[4347] = 1'd0;
    assign memhint[4348] = 1'd0;
    assign memhint[4349] = 1'd0;
    assign memhint[4350] = 1'd0;
    assign memhint[4351] = 1'd0;
    assign memhint[4352] = 1'd0;
    assign memhint[4353] = 1'd0;
    assign memhint[4354] = 1'd0;
    assign memhint[4355] = 1'd0;
    assign memhint[4356] = 1'd0;
    assign memhint[4357] = 1'd1;
    assign memhint[4358] = 1'd1;
    assign memhint[4359] = 1'd0;
    assign memhint[4360] = 1'd0;
    assign memhint[4361] = 1'd0;
    assign memhint[4362] = 1'd0;
    assign memhint[4363] = 1'd0;
    assign memhint[4364] = 1'd0;
    assign memhint[4365] = 1'd0;
    assign memhint[4366] = 1'd0;
    assign memhint[4367] = 1'd1;
    assign memhint[4368] = 1'd1;
    assign memhint[4369] = 1'd0;
    assign memhint[4370] = 1'd0;
    assign memhint[4371] = 1'd0;
    assign memhint[4372] = 1'd0;
    assign memhint[4373] = 1'd0;
    assign memhint[4374] = 1'd0;
    assign memhint[4375] = 1'd0;
    assign memhint[4376] = 1'd0;
    assign memhint[4377] = 1'd0;
    assign memhint[4378] = 1'd0;
    assign memhint[4379] = 1'd0;
    assign memhint[4380] = 1'd0;
    assign memhint[4381] = 1'd0;
    assign memhint[4382] = 1'd0;
    assign memhint[4383] = 1'd0;
    assign memhint[4384] = 1'd0;
    assign memhint[4385] = 1'd0;
    assign memhint[4386] = 1'd0;
    assign memhint[4387] = 1'd0;
    assign memhint[4388] = 1'd0;
    assign memhint[4389] = 1'd1;
    assign memhint[4390] = 1'd1;
    assign memhint[4391] = 1'd0;
    assign memhint[4392] = 1'd0;
    assign memhint[4393] = 1'd0;
    assign memhint[4394] = 1'd0;
    assign memhint[4395] = 1'd0;
    assign memhint[4396] = 1'd0;
    assign memhint[4397] = 1'd0;
    assign memhint[4398] = 1'd0;
    assign memhint[4399] = 1'd0;
    assign memhint[4400] = 1'd0;
    assign memhint[4401] = 1'd0;
    assign memhint[4402] = 1'd0;
    assign memhint[4403] = 1'd0;
    assign memhint[4404] = 1'd0;
    assign memhint[4405] = 1'd1;
    assign memhint[4406] = 1'd1;
    assign memhint[4407] = 1'd1;
    assign memhint[4408] = 1'd1;
    assign memhint[4409] = 1'd1;
    assign memhint[4410] = 1'd1;
    assign memhint[4411] = 1'd1;
    assign memhint[4412] = 1'd1;
    assign memhint[4413] = 1'd1;
    assign memhint[4414] = 1'd1;
    assign memhint[4415] = 1'd0;
    assign memhint[4416] = 1'd0;
    assign memhint[4417] = 1'd0;
    assign memhint[4418] = 1'd0;
    assign memhint[4419] = 1'd0;
    assign memhint[4420] = 1'd0;
    assign memhint[4421] = 1'd0;
    assign memhint[4422] = 1'd0;
    assign memhint[4423] = 1'd0;
    assign memhint[4424] = 1'd1;
    assign memhint[4425] = 1'd1;
    assign memhint[4426] = 1'd0;
    assign memhint[4427] = 1'd0;
    assign memhint[4428] = 1'd0;
    assign memhint[4429] = 1'd0;
    assign memhint[4430] = 1'd0;
    assign memhint[4431] = 1'd0;
    assign memhint[4432] = 1'd0;
    assign memhint[4433] = 1'd0;
    assign memhint[4434] = 1'd0;
    assign memhint[4435] = 1'd0;
    assign memhint[4436] = 1'd0;
    assign memhint[4437] = 1'd0;
    assign memhint[4438] = 1'd0;
    assign memhint[4439] = 1'd0;
    assign memhint[4440] = 1'd0;
    assign memhint[4441] = 1'd0;
    assign memhint[4442] = 1'd1;
    assign memhint[4443] = 1'd1;
    assign memhint[4444] = 1'd0;
    assign memhint[4445] = 1'd0;
    assign memhint[4446] = 1'd0;
    assign memhint[4447] = 1'd0;
    assign memhint[4448] = 1'd0;
    assign memhint[4449] = 1'd0;
    assign memhint[4450] = 1'd0;
    assign memhint[4451] = 1'd1;
    assign memhint[4452] = 1'd1;
    assign memhint[4453] = 1'd0;
    assign memhint[4454] = 1'd0;
    assign memhint[4455] = 1'd0;
    assign memhint[4456] = 1'd0;
    assign memhint[4457] = 1'd0;
    assign memhint[4458] = 1'd0;
    assign memhint[4459] = 1'd0;
    assign memhint[4460] = 1'd0;
    assign memhint[4461] = 1'd0;
    assign memhint[4462] = 1'd0;
    assign memhint[4463] = 1'd0;
    assign memhint[4464] = 1'd0;
    assign memhint[4465] = 1'd0;
    assign memhint[4466] = 1'd0;
    assign memhint[4467] = 1'd1;
    assign memhint[4468] = 1'd1;
    assign memhint[4469] = 1'd0;
    assign memhint[4470] = 1'd0;
    assign memhint[4471] = 1'd0;
    assign memhint[4472] = 1'd0;
    assign memhint[4473] = 1'd0;
    assign memhint[4474] = 1'd0;
    assign memhint[4475] = 1'd0;
    assign memhint[4476] = 1'd0;
    assign memhint[4477] = 1'd0;
    assign memhint[4478] = 1'd0;
    assign memhint[4479] = 1'd0;
    assign memhint[4480] = 1'd0;
    assign memhint[4481] = 1'd0;
    assign memhint[4482] = 1'd0;
    assign memhint[4483] = 1'd1;
    assign memhint[4484] = 1'd1;
    assign memhint[4485] = 1'd1;
    assign memhint[4486] = 1'd1;
    assign memhint[4487] = 1'd0;
    assign memhint[4488] = 1'd0;
    assign memhint[4489] = 1'd0;
    assign memhint[4490] = 1'd0;
    assign memhint[4491] = 1'd0;
    assign memhint[4492] = 1'd0;
    assign memhint[4493] = 1'd0;
    assign memhint[4494] = 1'd1;
    assign memhint[4495] = 1'd1;
    assign memhint[4496] = 1'd0;
    assign memhint[4497] = 1'd0;
    assign memhint[4498] = 1'd0;
    assign memhint[4499] = 1'd0;
    assign memhint[4500] = 1'd0;
    assign memhint[4501] = 1'd0;
    assign memhint[4502] = 1'd0;
    assign memhint[4503] = 1'd0;
    assign memhint[4504] = 1'd0;
    assign memhint[4505] = 1'd0;
    assign memhint[4506] = 1'd0;
    assign memhint[4507] = 1'd0;
    assign memhint[4508] = 1'd0;
    assign memhint[4509] = 1'd0;
    assign memhint[4510] = 1'd0;
    assign memhint[4511] = 1'd1;
    assign memhint[4512] = 1'd1;
    assign memhint[4513] = 1'd0;
    assign memhint[4514] = 1'd0;
    assign memhint[4515] = 1'd0;
    assign memhint[4516] = 1'd0;
    assign memhint[4517] = 1'd0;
    assign memhint[4518] = 1'd0;
    assign memhint[4519] = 1'd0;
    assign memhint[4520] = 1'd0;
    assign memhint[4521] = 1'd0;
    assign memhint[4522] = 1'd0;
    assign memhint[4523] = 1'd0;
    assign memhint[4524] = 1'd0;
    assign memhint[4525] = 1'd0;
    assign memhint[4526] = 1'd1;
    assign memhint[4527] = 1'd1;
    assign memhint[4528] = 1'd0;
    assign memhint[4529] = 1'd0;
    assign memhint[4530] = 1'd0;
    assign memhint[4531] = 1'd0;
    assign memhint[4532] = 1'd0;
    assign memhint[4533] = 1'd0;
    assign memhint[4534] = 1'd0;
    assign memhint[4535] = 1'd0;
    assign memhint[4536] = 1'd0;
    assign memhint[4537] = 1'd0;
    assign memhint[4538] = 1'd0;
    assign memhint[4539] = 1'd0;
    assign memhint[4540] = 1'd0;
    assign memhint[4541] = 1'd0;
    assign memhint[4542] = 1'd1;
    assign memhint[4543] = 1'd1;
    assign memhint[4544] = 1'd0;
    assign memhint[4545] = 1'd0;
    assign memhint[4546] = 1'd0;
    assign memhint[4547] = 1'd0;
    assign memhint[4548] = 1'd0;
    assign memhint[4549] = 1'd0;
    assign memhint[4550] = 1'd0;
    assign memhint[4551] = 1'd0;
    assign memhint[4552] = 1'd0;
    assign memhint[4553] = 1'd0;
    assign memhint[4554] = 1'd0;
    assign memhint[4555] = 1'd0;
    assign memhint[4556] = 1'd0;
    assign memhint[4557] = 1'd0;
    assign memhint[4558] = 1'd0;
    assign memhint[4559] = 1'd0;
    assign memhint[4560] = 1'd0;
    assign memhint[4561] = 1'd0;
    assign memhint[4562] = 1'd0;
    assign memhint[4563] = 1'd0;
    assign memhint[4564] = 1'd0;
    assign memhint[4565] = 1'd0;
    assign memhint[4566] = 1'd0;
    assign memhint[4567] = 1'd0;
    assign memhint[4568] = 1'd0;
    assign memhint[4569] = 1'd0;
    assign memhint[4570] = 1'd0;
    assign memhint[4571] = 1'd1;
    assign memhint[4572] = 1'd1;
    assign memhint[4573] = 1'd0;
    assign memhint[4574] = 1'd0;
    assign memhint[4575] = 1'd0;
    assign memhint[4576] = 1'd0;
    assign memhint[4577] = 1'd0;
    assign memhint[4578] = 1'd0;
    assign memhint[4579] = 1'd0;
    assign memhint[4580] = 1'd0;
    assign memhint[4581] = 1'd0;
    assign memhint[4582] = 1'd0;
    assign memhint[4583] = 1'd0;
    assign memhint[4584] = 1'd0;
    assign memhint[4585] = 1'd0;
    assign memhint[4586] = 1'd0;
    assign memhint[4587] = 1'd0;
    assign memhint[4588] = 1'd0;
    assign memhint[4589] = 1'd0;
    assign memhint[4590] = 1'd0;
    assign memhint[4591] = 1'd0;
    assign memhint[4592] = 1'd0;
    assign memhint[4593] = 1'd0;
    assign memhint[4594] = 1'd1;
    assign memhint[4595] = 1'd1;
    assign memhint[4596] = 1'd0;
    assign memhint[4597] = 1'd0;
    assign memhint[4598] = 1'd0;
    assign memhint[4599] = 1'd0;
    assign memhint[4600] = 1'd0;
    assign memhint[4601] = 1'd0;
    assign memhint[4602] = 1'd0;
    assign memhint[4603] = 1'd1;
    assign memhint[4604] = 1'd1;
    assign memhint[4605] = 1'd0;
    assign memhint[4606] = 1'd0;
    assign memhint[4607] = 1'd0;
    assign memhint[4608] = 1'd0;
    assign memhint[4609] = 1'd0;
    assign memhint[4610] = 1'd0;
    assign memhint[4611] = 1'd0;
    assign memhint[4612] = 1'd0;
    assign memhint[4613] = 1'd0;
    assign memhint[4614] = 1'd0;
    assign memhint[4615] = 1'd0;
    assign memhint[4616] = 1'd0;
    assign memhint[4617] = 1'd0;
    assign memhint[4618] = 1'd0;
    assign memhint[4619] = 1'd0;
    assign memhint[4620] = 1'd0;
    assign memhint[4621] = 1'd0;
    assign memhint[4622] = 1'd0;
    assign memhint[4623] = 1'd0;
    assign memhint[4624] = 1'd0;
    assign memhint[4625] = 1'd0;
    assign memhint[4626] = 1'd0;
    assign memhint[4627] = 1'd0;
    assign memhint[4628] = 1'd1;
    assign memhint[4629] = 1'd1;
    assign memhint[4630] = 1'd1;
    assign memhint[4631] = 1'd1;
    assign memhint[4632] = 1'd0;
    assign memhint[4633] = 1'd0;
    assign memhint[4634] = 1'd0;
    assign memhint[4635] = 1'd0;
    assign memhint[4636] = 1'd0;
    assign memhint[4637] = 1'd0;
    assign memhint[4638] = 1'd1;
    assign memhint[4639] = 1'd1;
    assign memhint[4640] = 1'd0;
    assign memhint[4641] = 1'd0;
    assign memhint[4642] = 1'd0;
    assign memhint[4643] = 1'd0;
    assign memhint[4644] = 1'd0;
    assign memhint[4645] = 1'd0;
    assign memhint[4646] = 1'd0;
    assign memhint[4647] = 1'd0;
    assign memhint[4648] = 1'd0;
    assign memhint[4649] = 1'd0;
    assign memhint[4650] = 1'd0;
    assign memhint[4651] = 1'd0;
    assign memhint[4652] = 1'd0;
    assign memhint[4653] = 1'd0;
    assign memhint[4654] = 1'd0;
    assign memhint[4655] = 1'd0;
    assign memhint[4656] = 1'd0;
    assign memhint[4657] = 1'd0;
    assign memhint[4658] = 1'd0;
    assign memhint[4659] = 1'd0;
    assign memhint[4660] = 1'd1;
    assign memhint[4661] = 1'd1;
    assign memhint[4662] = 1'd0;
    assign memhint[4663] = 1'd0;
    assign memhint[4664] = 1'd0;
    assign memhint[4665] = 1'd0;
    assign memhint[4666] = 1'd0;
    assign memhint[4667] = 1'd1;
    assign memhint[4668] = 1'd1;
    assign memhint[4669] = 1'd0;
    assign memhint[4670] = 1'd0;
    assign memhint[4671] = 1'd0;
    assign memhint[4672] = 1'd0;
    assign memhint[4673] = 1'd0;
    assign memhint[4674] = 1'd0;
    assign memhint[4675] = 1'd0;
    assign memhint[4676] = 1'd1;
    assign memhint[4677] = 1'd1;
    assign memhint[4678] = 1'd0;
    assign memhint[4679] = 1'd0;
    assign memhint[4680] = 1'd0;
    assign memhint[4681] = 1'd0;
    assign memhint[4682] = 1'd0;
    assign memhint[4683] = 1'd1;
    assign memhint[4684] = 1'd1;
    assign memhint[4685] = 1'd0;
    assign memhint[4686] = 1'd0;
    assign memhint[4687] = 1'd0;
    assign memhint[4688] = 1'd0;
    assign memhint[4689] = 1'd0;
    assign memhint[4690] = 1'd1;
    assign memhint[4691] = 1'd1;
    assign memhint[4692] = 1'd0;
    assign memhint[4693] = 1'd0;
    assign memhint[4694] = 1'd0;
    assign memhint[4695] = 1'd0;
    assign memhint[4696] = 1'd0;
    assign memhint[4697] = 1'd0;
    assign memhint[4698] = 1'd0;
    assign memhint[4699] = 1'd0;
    assign memhint[4700] = 1'd0;
    assign memhint[4701] = 1'd0;
    assign memhint[4702] = 1'd0;
    assign memhint[4703] = 1'd0;
    assign memhint[4704] = 1'd1;
    assign memhint[4705] = 1'd1;
    assign memhint[4706] = 1'd1;
    assign memhint[4707] = 1'd1;
    assign memhint[4708] = 1'd1;
    assign memhint[4709] = 1'd1;
    assign memhint[4710] = 1'd1;
    assign memhint[4711] = 1'd1;
    assign memhint[4712] = 1'd1;
    assign memhint[4713] = 1'd1;
    assign memhint[4714] = 1'd0;
    assign memhint[4715] = 1'd0;
    assign memhint[4716] = 1'd0;
    assign memhint[4717] = 1'd0;
    assign memhint[4718] = 1'd0;
    assign memhint[4719] = 1'd0;
    assign memhint[4720] = 1'd0;
    assign memhint[4721] = 1'd0;
    assign memhint[4722] = 1'd0;
    assign memhint[4723] = 1'd0;
    assign memhint[4724] = 1'd0;
    assign memhint[4725] = 1'd0;
    assign memhint[4726] = 1'd0;
    assign memhint[4727] = 1'd0;
    assign memhint[4728] = 1'd0;
    assign memhint[4729] = 1'd0;
    assign memhint[4730] = 1'd1;
    assign memhint[4731] = 1'd1;
    assign memhint[4732] = 1'd0;
    assign memhint[4733] = 1'd0;
    assign memhint[4734] = 1'd0;
    assign memhint[4735] = 1'd0;
    assign memhint[4736] = 1'd0;
    assign memhint[4737] = 1'd0;
    assign memhint[4738] = 1'd0;
    assign memhint[4739] = 1'd0;
    assign memhint[4740] = 1'd1;
    assign memhint[4741] = 1'd1;
    assign memhint[4742] = 1'd0;
    assign memhint[4743] = 1'd0;
    assign memhint[4744] = 1'd0;
    assign memhint[4745] = 1'd0;
    assign memhint[4746] = 1'd0;
    assign memhint[4747] = 1'd0;
    assign memhint[4748] = 1'd0;
    assign memhint[4749] = 1'd0;
    assign memhint[4750] = 1'd0;
    assign memhint[4751] = 1'd0;
    assign memhint[4752] = 1'd0;
    assign memhint[4753] = 1'd0;
    assign memhint[4754] = 1'd0;
    assign memhint[4755] = 1'd0;
    assign memhint[4756] = 1'd0;
    assign memhint[4757] = 1'd0;
    assign memhint[4758] = 1'd0;
    assign memhint[4759] = 1'd0;
    assign memhint[4760] = 1'd0;
    assign memhint[4761] = 1'd0;
    assign memhint[4762] = 1'd1;
    assign memhint[4763] = 1'd1;
    assign memhint[4764] = 1'd0;
    assign memhint[4765] = 1'd0;
    assign memhint[4766] = 1'd0;
    assign memhint[4767] = 1'd0;
    assign memhint[4768] = 1'd0;
    assign memhint[4769] = 1'd0;
    assign memhint[4770] = 1'd0;
    assign memhint[4771] = 1'd0;
    assign memhint[4772] = 1'd0;
    assign memhint[4773] = 1'd0;
    assign memhint[4774] = 1'd0;
    assign memhint[4775] = 1'd0;
    assign memhint[4776] = 1'd0;
    assign memhint[4777] = 1'd0;
    assign memhint[4778] = 1'd1;
    assign memhint[4779] = 1'd1;
    assign memhint[4780] = 1'd0;
    assign memhint[4781] = 1'd0;
    assign memhint[4782] = 1'd0;
    assign memhint[4783] = 1'd0;
    assign memhint[4784] = 1'd0;
    assign memhint[4785] = 1'd0;
    assign memhint[4786] = 1'd0;
    assign memhint[4787] = 1'd0;
    assign memhint[4788] = 1'd0;
    assign memhint[4789] = 1'd0;
    assign memhint[4790] = 1'd0;
    assign memhint[4791] = 1'd0;
    assign memhint[4792] = 1'd0;
    assign memhint[4793] = 1'd0;
    assign memhint[4794] = 1'd0;
    assign memhint[4795] = 1'd0;
    assign memhint[4796] = 1'd0;
    assign memhint[4797] = 1'd1;
    assign memhint[4798] = 1'd1;
    assign memhint[4799] = 1'd0;
    assign memhint[4800] = 1'd0;
    assign memhint[4801] = 1'd0;
    assign memhint[4802] = 1'd0;
    assign memhint[4803] = 1'd0;
    assign memhint[4804] = 1'd0;
    assign memhint[4805] = 1'd0;
    assign memhint[4806] = 1'd0;
    assign memhint[4807] = 1'd0;
    assign memhint[4808] = 1'd0;
    assign memhint[4809] = 1'd0;
    assign memhint[4810] = 1'd0;
    assign memhint[4811] = 1'd0;
    assign memhint[4812] = 1'd0;
    assign memhint[4813] = 1'd0;
    assign memhint[4814] = 1'd0;
    assign memhint[4815] = 1'd1;
    assign memhint[4816] = 1'd1;
    assign memhint[4817] = 1'd0;
    assign memhint[4818] = 1'd0;
    assign memhint[4819] = 1'd0;
    assign memhint[4820] = 1'd0;
    assign memhint[4821] = 1'd0;
    assign memhint[4822] = 1'd0;
    assign memhint[4823] = 1'd0;
    assign memhint[4824] = 1'd1;
    assign memhint[4825] = 1'd1;
    assign memhint[4826] = 1'd0;
    assign memhint[4827] = 1'd0;
    assign memhint[4828] = 1'd0;
    assign memhint[4829] = 1'd0;
    assign memhint[4830] = 1'd0;
    assign memhint[4831] = 1'd0;
    assign memhint[4832] = 1'd0;
    assign memhint[4833] = 1'd0;
    assign memhint[4834] = 1'd0;
    assign memhint[4835] = 1'd0;
    assign memhint[4836] = 1'd0;
    assign memhint[4837] = 1'd0;
    assign memhint[4838] = 1'd0;
    assign memhint[4839] = 1'd0;
    assign memhint[4840] = 1'd1;
    assign memhint[4841] = 1'd1;
    assign memhint[4842] = 1'd0;
    assign memhint[4843] = 1'd0;
    assign memhint[4844] = 1'd0;
    assign memhint[4845] = 1'd0;
    assign memhint[4846] = 1'd0;
    assign memhint[4847] = 1'd0;
    assign memhint[4848] = 1'd0;
    assign memhint[4849] = 1'd0;
    assign memhint[4850] = 1'd0;
    assign memhint[4851] = 1'd0;
    assign memhint[4852] = 1'd0;
    assign memhint[4853] = 1'd0;
    assign memhint[4854] = 1'd0;
    assign memhint[4855] = 1'd0;
    assign memhint[4856] = 1'd0;
    assign memhint[4857] = 1'd0;
    assign memhint[4858] = 1'd1;
    assign memhint[4859] = 1'd1;
    assign memhint[4860] = 1'd1;
    assign memhint[4861] = 1'd0;
    assign memhint[4862] = 1'd0;
    assign memhint[4863] = 1'd0;
    assign memhint[4864] = 1'd0;
    assign memhint[4865] = 1'd0;
    assign memhint[4866] = 1'd0;
    assign memhint[4867] = 1'd1;
    assign memhint[4868] = 1'd1;
    assign memhint[4869] = 1'd0;
    assign memhint[4870] = 1'd0;
    assign memhint[4871] = 1'd0;
    assign memhint[4872] = 1'd0;
    assign memhint[4873] = 1'd0;
    assign memhint[4874] = 1'd0;
    assign memhint[4875] = 1'd0;
    assign memhint[4876] = 1'd0;
    assign memhint[4877] = 1'd0;
    assign memhint[4878] = 1'd0;
    assign memhint[4879] = 1'd0;
    assign memhint[4880] = 1'd0;
    assign memhint[4881] = 1'd0;
    assign memhint[4882] = 1'd0;
    assign memhint[4883] = 1'd0;
    assign memhint[4884] = 1'd1;
    assign memhint[4885] = 1'd1;
    assign memhint[4886] = 1'd0;
    assign memhint[4887] = 1'd0;
    assign memhint[4888] = 1'd0;
    assign memhint[4889] = 1'd0;
    assign memhint[4890] = 1'd0;
    assign memhint[4891] = 1'd0;
    assign memhint[4892] = 1'd0;
    assign memhint[4893] = 1'd0;
    assign memhint[4894] = 1'd0;
    assign memhint[4895] = 1'd0;
    assign memhint[4896] = 1'd0;
    assign memhint[4897] = 1'd0;
    assign memhint[4898] = 1'd0;
    assign memhint[4899] = 1'd1;
    assign memhint[4900] = 1'd1;
    assign memhint[4901] = 1'd0;
    assign memhint[4902] = 1'd0;
    assign memhint[4903] = 1'd0;
    assign memhint[4904] = 1'd0;
    assign memhint[4905] = 1'd0;
    assign memhint[4906] = 1'd0;
    assign memhint[4907] = 1'd0;
    assign memhint[4908] = 1'd0;
    assign memhint[4909] = 1'd0;
    assign memhint[4910] = 1'd0;
    assign memhint[4911] = 1'd0;
    assign memhint[4912] = 1'd0;
    assign memhint[4913] = 1'd0;
    assign memhint[4914] = 1'd0;
    assign memhint[4915] = 1'd1;
    assign memhint[4916] = 1'd1;
    assign memhint[4917] = 1'd0;
    assign memhint[4918] = 1'd0;
    assign memhint[4919] = 1'd0;
    assign memhint[4920] = 1'd0;
    assign memhint[4921] = 1'd0;
    assign memhint[4922] = 1'd0;
    assign memhint[4923] = 1'd0;
    assign memhint[4924] = 1'd0;
    assign memhint[4925] = 1'd0;
    assign memhint[4926] = 1'd0;
    assign memhint[4927] = 1'd0;
    assign memhint[4928] = 1'd0;
    assign memhint[4929] = 1'd0;
    assign memhint[4930] = 1'd0;
    assign memhint[4931] = 1'd0;
    assign memhint[4932] = 1'd0;
    assign memhint[4933] = 1'd0;
    assign memhint[4934] = 1'd0;
    assign memhint[4935] = 1'd0;
    assign memhint[4936] = 1'd0;
    assign memhint[4937] = 1'd0;
    assign memhint[4938] = 1'd0;
    assign memhint[4939] = 1'd0;
    assign memhint[4940] = 1'd0;
    assign memhint[4941] = 1'd0;
    assign memhint[4942] = 1'd0;
    assign memhint[4943] = 1'd0;
    assign memhint[4944] = 1'd1;
    assign memhint[4945] = 1'd1;
    assign memhint[4946] = 1'd0;
    assign memhint[4947] = 1'd0;
    assign memhint[4948] = 1'd0;
    assign memhint[4949] = 1'd0;
    assign memhint[4950] = 1'd0;
    assign memhint[4951] = 1'd0;
    assign memhint[4952] = 1'd0;
    assign memhint[4953] = 1'd0;
    assign memhint[4954] = 1'd0;
    assign memhint[4955] = 1'd0;
    assign memhint[4956] = 1'd0;
    assign memhint[4957] = 1'd0;
    assign memhint[4958] = 1'd0;
    assign memhint[4959] = 1'd0;
    assign memhint[4960] = 1'd0;
    assign memhint[4961] = 1'd0;
    assign memhint[4962] = 1'd0;
    assign memhint[4963] = 1'd0;
    assign memhint[4964] = 1'd0;
    assign memhint[4965] = 1'd0;
    assign memhint[4966] = 1'd1;
    assign memhint[4967] = 1'd1;
    assign memhint[4968] = 1'd1;
    assign memhint[4969] = 1'd1;
    assign memhint[4970] = 1'd1;
    assign memhint[4971] = 1'd1;
    assign memhint[4972] = 1'd1;
    assign memhint[4973] = 1'd1;
    assign memhint[4974] = 1'd1;
    assign memhint[4975] = 1'd1;
    assign memhint[4976] = 1'd1;
    assign memhint[4977] = 1'd1;
    assign memhint[4978] = 1'd1;
    assign memhint[4979] = 1'd0;
    assign memhint[4980] = 1'd0;
    assign memhint[4981] = 1'd0;
    assign memhint[4982] = 1'd0;
    assign memhint[4983] = 1'd0;
    assign memhint[4984] = 1'd0;
    assign memhint[4985] = 1'd0;
    assign memhint[4986] = 1'd0;
    assign memhint[4987] = 1'd0;
    assign memhint[4988] = 1'd0;
    assign memhint[4989] = 1'd0;
    assign memhint[4990] = 1'd0;
    assign memhint[4991] = 1'd0;
    assign memhint[4992] = 1'd0;
    assign memhint[4993] = 1'd0;
    assign memhint[4994] = 1'd0;
    assign memhint[4995] = 1'd0;
    assign memhint[4996] = 1'd0;
    assign memhint[4997] = 1'd0;
    assign memhint[4998] = 1'd0;
    assign memhint[4999] = 1'd0;
    assign memhint[5000] = 1'd0;
    assign memhint[5001] = 1'd0;
    assign memhint[5002] = 1'd0;
    assign memhint[5003] = 1'd1;
    assign memhint[5004] = 1'd1;
    assign memhint[5005] = 1'd1;
    assign memhint[5006] = 1'd0;
    assign memhint[5007] = 1'd0;
    assign memhint[5008] = 1'd0;
    assign memhint[5009] = 1'd0;
    assign memhint[5010] = 1'd0;
    assign memhint[5011] = 1'd1;
    assign memhint[5012] = 1'd1;
    assign memhint[5013] = 1'd0;
    assign memhint[5014] = 1'd0;
    assign memhint[5015] = 1'd0;
    assign memhint[5016] = 1'd0;
    assign memhint[5017] = 1'd0;
    assign memhint[5018] = 1'd0;
    assign memhint[5019] = 1'd0;
    assign memhint[5020] = 1'd0;
    assign memhint[5021] = 1'd0;
    assign memhint[5022] = 1'd0;
    assign memhint[5023] = 1'd0;
    assign memhint[5024] = 1'd0;
    assign memhint[5025] = 1'd0;
    assign memhint[5026] = 1'd0;
    assign memhint[5027] = 1'd0;
    assign memhint[5028] = 1'd0;
    assign memhint[5029] = 1'd0;
    assign memhint[5030] = 1'd0;
    assign memhint[5031] = 1'd0;
    assign memhint[5032] = 1'd0;
    assign memhint[5033] = 1'd1;
    assign memhint[5034] = 1'd1;
    assign memhint[5035] = 1'd0;
    assign memhint[5036] = 1'd0;
    assign memhint[5037] = 1'd0;
    assign memhint[5038] = 1'd0;
    assign memhint[5039] = 1'd0;
    assign memhint[5040] = 1'd1;
    assign memhint[5041] = 1'd1;
    assign memhint[5042] = 1'd0;
    assign memhint[5043] = 1'd0;
    assign memhint[5044] = 1'd0;
    assign memhint[5045] = 1'd0;
    assign memhint[5046] = 1'd0;
    assign memhint[5047] = 1'd0;
    assign memhint[5048] = 1'd0;
    assign memhint[5049] = 1'd0;
    assign memhint[5050] = 1'd1;
    assign memhint[5051] = 1'd1;
    assign memhint[5052] = 1'd0;
    assign memhint[5053] = 1'd0;
    assign memhint[5054] = 1'd0;
    assign memhint[5055] = 1'd0;
    assign memhint[5056] = 1'd1;
    assign memhint[5057] = 1'd1;
    assign memhint[5058] = 1'd0;
    assign memhint[5059] = 1'd0;
    assign memhint[5060] = 1'd0;
    assign memhint[5061] = 1'd0;
    assign memhint[5062] = 1'd0;
    assign memhint[5063] = 1'd1;
    assign memhint[5064] = 1'd1;
    assign memhint[5065] = 1'd0;
    assign memhint[5066] = 1'd0;
    assign memhint[5067] = 1'd0;
    assign memhint[5068] = 1'd0;
    assign memhint[5069] = 1'd0;
    assign memhint[5070] = 1'd0;
    assign memhint[5071] = 1'd0;
    assign memhint[5072] = 1'd0;
    assign memhint[5073] = 1'd0;
    assign memhint[5074] = 1'd0;
    assign memhint[5075] = 1'd0;
    assign memhint[5076] = 1'd0;
    assign memhint[5077] = 1'd1;
    assign memhint[5078] = 1'd1;
    assign memhint[5079] = 1'd1;
    assign memhint[5080] = 1'd1;
    assign memhint[5081] = 1'd1;
    assign memhint[5082] = 1'd1;
    assign memhint[5083] = 1'd1;
    assign memhint[5084] = 1'd1;
    assign memhint[5085] = 1'd1;
    assign memhint[5086] = 1'd1;
    assign memhint[5087] = 1'd0;
    assign memhint[5088] = 1'd0;
    assign memhint[5089] = 1'd0;
    assign memhint[5090] = 1'd0;
    assign memhint[5091] = 1'd0;
    assign memhint[5092] = 1'd0;
    assign memhint[5093] = 1'd0;
    assign memhint[5094] = 1'd0;
    assign memhint[5095] = 1'd0;
    assign memhint[5096] = 1'd0;
    assign memhint[5097] = 1'd0;
    assign memhint[5098] = 1'd0;
    assign memhint[5099] = 1'd0;
    assign memhint[5100] = 1'd0;
    assign memhint[5101] = 1'd0;
    assign memhint[5102] = 1'd0;
    assign memhint[5103] = 1'd1;
    assign memhint[5104] = 1'd1;
    assign memhint[5105] = 1'd0;
    assign memhint[5106] = 1'd0;
    assign memhint[5107] = 1'd0;
    assign memhint[5108] = 1'd0;
    assign memhint[5109] = 1'd0;
    assign memhint[5110] = 1'd0;
    assign memhint[5111] = 1'd0;
    assign memhint[5112] = 1'd0;
    assign memhint[5113] = 1'd1;
    assign memhint[5114] = 1'd1;
    assign memhint[5115] = 1'd0;
    assign memhint[5116] = 1'd0;
    assign memhint[5117] = 1'd0;
    assign memhint[5118] = 1'd0;
    assign memhint[5119] = 1'd0;
    assign memhint[5120] = 1'd0;
    assign memhint[5121] = 1'd0;
    assign memhint[5122] = 1'd0;
    assign memhint[5123] = 1'd0;
    assign memhint[5124] = 1'd0;
    assign memhint[5125] = 1'd0;
    assign memhint[5126] = 1'd0;
    assign memhint[5127] = 1'd0;
    assign memhint[5128] = 1'd0;
    assign memhint[5129] = 1'd0;
    assign memhint[5130] = 1'd0;
    assign memhint[5131] = 1'd0;
    assign memhint[5132] = 1'd0;
    assign memhint[5133] = 1'd0;
    assign memhint[5134] = 1'd0;
    assign memhint[5135] = 1'd1;
    assign memhint[5136] = 1'd1;
    assign memhint[5137] = 1'd0;
    assign memhint[5138] = 1'd0;
    assign memhint[5139] = 1'd0;
    assign memhint[5140] = 1'd0;
    assign memhint[5141] = 1'd0;
    assign memhint[5142] = 1'd0;
    assign memhint[5143] = 1'd0;
    assign memhint[5144] = 1'd0;
    assign memhint[5145] = 1'd0;
    assign memhint[5146] = 1'd0;
    assign memhint[5147] = 1'd0;
    assign memhint[5148] = 1'd0;
    assign memhint[5149] = 1'd0;
    assign memhint[5150] = 1'd0;
    assign memhint[5151] = 1'd1;
    assign memhint[5152] = 1'd1;
    assign memhint[5153] = 1'd0;
    assign memhint[5154] = 1'd0;
    assign memhint[5155] = 1'd0;
    assign memhint[5156] = 1'd0;
    assign memhint[5157] = 1'd0;
    assign memhint[5158] = 1'd0;
    assign memhint[5159] = 1'd0;
    assign memhint[5160] = 1'd0;
    assign memhint[5161] = 1'd0;
    assign memhint[5162] = 1'd0;
    assign memhint[5163] = 1'd0;
    assign memhint[5164] = 1'd0;
    assign memhint[5165] = 1'd0;
    assign memhint[5166] = 1'd0;
    assign memhint[5167] = 1'd0;
    assign memhint[5168] = 1'd0;
    assign memhint[5169] = 1'd0;
    assign memhint[5170] = 1'd1;
    assign memhint[5171] = 1'd1;
    assign memhint[5172] = 1'd0;
    assign memhint[5173] = 1'd0;
    assign memhint[5174] = 1'd0;
    assign memhint[5175] = 1'd0;
    assign memhint[5176] = 1'd0;
    assign memhint[5177] = 1'd0;
    assign memhint[5178] = 1'd0;
    assign memhint[5179] = 1'd0;
    assign memhint[5180] = 1'd0;
    assign memhint[5181] = 1'd0;
    assign memhint[5182] = 1'd0;
    assign memhint[5183] = 1'd0;
    assign memhint[5184] = 1'd0;
    assign memhint[5185] = 1'd0;
    assign memhint[5186] = 1'd0;
    assign memhint[5187] = 1'd1;
    assign memhint[5188] = 1'd1;
    assign memhint[5189] = 1'd1;
    assign memhint[5190] = 1'd1;
    assign memhint[5191] = 1'd1;
    assign memhint[5192] = 1'd1;
    assign memhint[5193] = 1'd1;
    assign memhint[5194] = 1'd1;
    assign memhint[5195] = 1'd1;
    assign memhint[5196] = 1'd1;
    assign memhint[5197] = 1'd1;
    assign memhint[5198] = 1'd1;
    assign memhint[5199] = 1'd1;
    assign memhint[5200] = 1'd0;
    assign memhint[5201] = 1'd0;
    assign memhint[5202] = 1'd0;
    assign memhint[5203] = 1'd0;
    assign memhint[5204] = 1'd0;
    assign memhint[5205] = 1'd0;
    assign memhint[5206] = 1'd0;
    assign memhint[5207] = 1'd0;
    assign memhint[5208] = 1'd0;
    assign memhint[5209] = 1'd0;
    assign memhint[5210] = 1'd0;
    assign memhint[5211] = 1'd0;
    assign memhint[5212] = 1'd0;
    assign memhint[5213] = 1'd1;
    assign memhint[5214] = 1'd1;
    assign memhint[5215] = 1'd0;
    assign memhint[5216] = 1'd0;
    assign memhint[5217] = 1'd0;
    assign memhint[5218] = 1'd0;
    assign memhint[5219] = 1'd0;
    assign memhint[5220] = 1'd0;
    assign memhint[5221] = 1'd0;
    assign memhint[5222] = 1'd0;
    assign memhint[5223] = 1'd0;
    assign memhint[5224] = 1'd0;
    assign memhint[5225] = 1'd0;
    assign memhint[5226] = 1'd0;
    assign memhint[5227] = 1'd0;
    assign memhint[5228] = 1'd0;
    assign memhint[5229] = 1'd0;
    assign memhint[5230] = 1'd0;
    assign memhint[5231] = 1'd0;
    assign memhint[5232] = 1'd1;
    assign memhint[5233] = 1'd1;
    assign memhint[5234] = 1'd0;
    assign memhint[5235] = 1'd0;
    assign memhint[5236] = 1'd0;
    assign memhint[5237] = 1'd0;
    assign memhint[5238] = 1'd0;
    assign memhint[5239] = 1'd0;
    assign memhint[5240] = 1'd1;
    assign memhint[5241] = 1'd1;
    assign memhint[5242] = 1'd0;
    assign memhint[5243] = 1'd0;
    assign memhint[5244] = 1'd0;
    assign memhint[5245] = 1'd0;
    assign memhint[5246] = 1'd0;
    assign memhint[5247] = 1'd0;
    assign memhint[5248] = 1'd0;
    assign memhint[5249] = 1'd0;
    assign memhint[5250] = 1'd0;
    assign memhint[5251] = 1'd0;
    assign memhint[5252] = 1'd0;
    assign memhint[5253] = 1'd0;
    assign memhint[5254] = 1'd0;
    assign memhint[5255] = 1'd0;
    assign memhint[5256] = 1'd0;
    assign memhint[5257] = 1'd1;
    assign memhint[5258] = 1'd1;
    assign memhint[5259] = 1'd0;
    assign memhint[5260] = 1'd0;
    assign memhint[5261] = 1'd0;
    assign memhint[5262] = 1'd0;
    assign memhint[5263] = 1'd0;
    assign memhint[5264] = 1'd0;
    assign memhint[5265] = 1'd0;
    assign memhint[5266] = 1'd0;
    assign memhint[5267] = 1'd0;
    assign memhint[5268] = 1'd0;
    assign memhint[5269] = 1'd0;
    assign memhint[5270] = 1'd0;
    assign memhint[5271] = 1'd0;
    assign memhint[5272] = 1'd1;
    assign memhint[5273] = 1'd1;
    assign memhint[5274] = 1'd0;
    assign memhint[5275] = 1'd0;
    assign memhint[5276] = 1'd0;
    assign memhint[5277] = 1'd0;
    assign memhint[5278] = 1'd0;
    assign memhint[5279] = 1'd0;
    assign memhint[5280] = 1'd0;
    assign memhint[5281] = 1'd0;
    assign memhint[5282] = 1'd0;
    assign memhint[5283] = 1'd0;
    assign memhint[5284] = 1'd0;
    assign memhint[5285] = 1'd0;
    assign memhint[5286] = 1'd0;
    assign memhint[5287] = 1'd0;
    assign memhint[5288] = 1'd1;
    assign memhint[5289] = 1'd1;
    assign memhint[5290] = 1'd0;
    assign memhint[5291] = 1'd0;
    assign memhint[5292] = 1'd0;
    assign memhint[5293] = 1'd0;
    assign memhint[5294] = 1'd0;
    assign memhint[5295] = 1'd0;
    assign memhint[5296] = 1'd0;
    assign memhint[5297] = 1'd0;
    assign memhint[5298] = 1'd0;
    assign memhint[5299] = 1'd0;
    assign memhint[5300] = 1'd0;
    assign memhint[5301] = 1'd0;
    assign memhint[5302] = 1'd0;
    assign memhint[5303] = 1'd0;
    assign memhint[5304] = 1'd0;
    assign memhint[5305] = 1'd0;
    assign memhint[5306] = 1'd0;
    assign memhint[5307] = 1'd0;
    assign memhint[5308] = 1'd0;
    assign memhint[5309] = 1'd0;
    assign memhint[5310] = 1'd0;
    assign memhint[5311] = 1'd0;
    assign memhint[5312] = 1'd0;
    assign memhint[5313] = 1'd0;
    assign memhint[5314] = 1'd0;
    assign memhint[5315] = 1'd0;
    assign memhint[5316] = 1'd0;
    assign memhint[5317] = 1'd1;
    assign memhint[5318] = 1'd1;
    assign memhint[5319] = 1'd0;
    assign memhint[5320] = 1'd0;
    assign memhint[5321] = 1'd0;
    assign memhint[5322] = 1'd0;
    assign memhint[5323] = 1'd0;
    assign memhint[5324] = 1'd0;
    assign memhint[5325] = 1'd0;
    assign memhint[5326] = 1'd0;
    assign memhint[5327] = 1'd0;
    assign memhint[5328] = 1'd0;
    assign memhint[5329] = 1'd0;
    assign memhint[5330] = 1'd0;
    assign memhint[5331] = 1'd0;
    assign memhint[5332] = 1'd0;
    assign memhint[5333] = 1'd0;
    assign memhint[5334] = 1'd0;
    assign memhint[5335] = 1'd0;
    assign memhint[5336] = 1'd0;
    assign memhint[5337] = 1'd0;
    assign memhint[5338] = 1'd0;
    assign memhint[5339] = 1'd1;
    assign memhint[5340] = 1'd1;
    assign memhint[5341] = 1'd1;
    assign memhint[5342] = 1'd1;
    assign memhint[5343] = 1'd1;
    assign memhint[5344] = 1'd1;
    assign memhint[5345] = 1'd1;
    assign memhint[5346] = 1'd1;
    assign memhint[5347] = 1'd1;
    assign memhint[5348] = 1'd1;
    assign memhint[5349] = 1'd1;
    assign memhint[5350] = 1'd1;
    assign memhint[5351] = 1'd1;
    assign memhint[5352] = 1'd0;
    assign memhint[5353] = 1'd0;
    assign memhint[5354] = 1'd0;
    assign memhint[5355] = 1'd0;
    assign memhint[5356] = 1'd0;
    assign memhint[5357] = 1'd0;
    assign memhint[5358] = 1'd0;
    assign memhint[5359] = 1'd0;
    assign memhint[5360] = 1'd0;
    assign memhint[5361] = 1'd0;
    assign memhint[5362] = 1'd0;
    assign memhint[5363] = 1'd0;
    assign memhint[5364] = 1'd0;
    assign memhint[5365] = 1'd0;
    assign memhint[5366] = 1'd0;
    assign memhint[5367] = 1'd0;
    assign memhint[5368] = 1'd0;
    assign memhint[5369] = 1'd0;
    assign memhint[5370] = 1'd0;
    assign memhint[5371] = 1'd0;
    assign memhint[5372] = 1'd0;
    assign memhint[5373] = 1'd0;
    assign memhint[5374] = 1'd0;
    assign memhint[5375] = 1'd0;
    assign memhint[5376] = 1'd0;
    assign memhint[5377] = 1'd1;
    assign memhint[5378] = 1'd1;
    assign memhint[5379] = 1'd0;
    assign memhint[5380] = 1'd0;
    assign memhint[5381] = 1'd0;
    assign memhint[5382] = 1'd0;
    assign memhint[5383] = 1'd0;
    assign memhint[5384] = 1'd1;
    assign memhint[5385] = 1'd1;
    assign memhint[5386] = 1'd0;
    assign memhint[5387] = 1'd0;
    assign memhint[5388] = 1'd0;
    assign memhint[5389] = 1'd0;
    assign memhint[5390] = 1'd0;
    assign memhint[5391] = 1'd0;
    assign memhint[5392] = 1'd0;
    assign memhint[5393] = 1'd0;
    assign memhint[5394] = 1'd0;
    assign memhint[5395] = 1'd0;
    assign memhint[5396] = 1'd0;
    assign memhint[5397] = 1'd0;
    assign memhint[5398] = 1'd0;
    assign memhint[5399] = 1'd0;
    assign memhint[5400] = 1'd0;
    assign memhint[5401] = 1'd0;
    assign memhint[5402] = 1'd0;
    assign memhint[5403] = 1'd0;
    assign memhint[5404] = 1'd0;
    assign memhint[5405] = 1'd0;
    assign memhint[5406] = 1'd1;
    assign memhint[5407] = 1'd1;
    assign memhint[5408] = 1'd0;
    assign memhint[5409] = 1'd0;
    assign memhint[5410] = 1'd0;
    assign memhint[5411] = 1'd0;
    assign memhint[5412] = 1'd0;
    assign memhint[5413] = 1'd1;
    assign memhint[5414] = 1'd1;
    assign memhint[5415] = 1'd0;
    assign memhint[5416] = 1'd0;
    assign memhint[5417] = 1'd0;
    assign memhint[5418] = 1'd0;
    assign memhint[5419] = 1'd0;
    assign memhint[5420] = 1'd0;
    assign memhint[5421] = 1'd0;
    assign memhint[5422] = 1'd0;
    assign memhint[5423] = 1'd1;
    assign memhint[5424] = 1'd1;
    assign memhint[5425] = 1'd1;
    assign memhint[5426] = 1'd0;
    assign memhint[5427] = 1'd0;
    assign memhint[5428] = 1'd0;
    assign memhint[5429] = 1'd1;
    assign memhint[5430] = 1'd1;
    assign memhint[5431] = 1'd0;
    assign memhint[5432] = 1'd0;
    assign memhint[5433] = 1'd0;
    assign memhint[5434] = 1'd0;
    assign memhint[5435] = 1'd0;
    assign memhint[5436] = 1'd1;
    assign memhint[5437] = 1'd1;
    assign memhint[5438] = 1'd1;
    assign memhint[5439] = 1'd0;
    assign memhint[5440] = 1'd0;
    assign memhint[5441] = 1'd0;
    assign memhint[5442] = 1'd0;
    assign memhint[5443] = 1'd0;
    assign memhint[5444] = 1'd0;
    assign memhint[5445] = 1'd0;
    assign memhint[5446] = 1'd0;
    assign memhint[5447] = 1'd0;
    assign memhint[5448] = 1'd0;
    assign memhint[5449] = 1'd0;
    assign memhint[5450] = 1'd0;
    assign memhint[5451] = 1'd0;
    assign memhint[5452] = 1'd0;
    assign memhint[5453] = 1'd0;
    assign memhint[5454] = 1'd0;
    assign memhint[5455] = 1'd0;
    assign memhint[5456] = 1'd0;
    assign memhint[5457] = 1'd0;
    assign memhint[5458] = 1'd1;
    assign memhint[5459] = 1'd1;
    assign memhint[5460] = 1'd0;
    assign memhint[5461] = 1'd0;
    assign memhint[5462] = 1'd0;
    assign memhint[5463] = 1'd0;
    assign memhint[5464] = 1'd0;
    assign memhint[5465] = 1'd0;
    assign memhint[5466] = 1'd0;
    assign memhint[5467] = 1'd0;
    assign memhint[5468] = 1'd0;
    assign memhint[5469] = 1'd0;
    assign memhint[5470] = 1'd0;
    assign memhint[5471] = 1'd0;
    assign memhint[5472] = 1'd0;
    assign memhint[5473] = 1'd0;
    assign memhint[5474] = 1'd0;
    assign memhint[5475] = 1'd0;
    assign memhint[5476] = 1'd1;
    assign memhint[5477] = 1'd1;
    assign memhint[5478] = 1'd0;
    assign memhint[5479] = 1'd0;
    assign memhint[5480] = 1'd0;
    assign memhint[5481] = 1'd0;
    assign memhint[5482] = 1'd0;
    assign memhint[5483] = 1'd0;
    assign memhint[5484] = 1'd0;
    assign memhint[5485] = 1'd0;
    assign memhint[5486] = 1'd1;
    assign memhint[5487] = 1'd1;
    assign memhint[5488] = 1'd0;
    assign memhint[5489] = 1'd0;
    assign memhint[5490] = 1'd0;
    assign memhint[5491] = 1'd0;
    assign memhint[5492] = 1'd0;
    assign memhint[5493] = 1'd0;
    assign memhint[5494] = 1'd0;
    assign memhint[5495] = 1'd0;
    assign memhint[5496] = 1'd0;
    assign memhint[5497] = 1'd0;
    assign memhint[5498] = 1'd0;
    assign memhint[5499] = 1'd0;
    assign memhint[5500] = 1'd0;
    assign memhint[5501] = 1'd0;
    assign memhint[5502] = 1'd0;
    assign memhint[5503] = 1'd0;
    assign memhint[5504] = 1'd0;
    assign memhint[5505] = 1'd0;
    assign memhint[5506] = 1'd0;
    assign memhint[5507] = 1'd0;
    assign memhint[5508] = 1'd1;
    assign memhint[5509] = 1'd1;
    assign memhint[5510] = 1'd0;
    assign memhint[5511] = 1'd0;
    assign memhint[5512] = 1'd0;
    assign memhint[5513] = 1'd0;
    assign memhint[5514] = 1'd0;
    assign memhint[5515] = 1'd0;
    assign memhint[5516] = 1'd0;
    assign memhint[5517] = 1'd0;
    assign memhint[5518] = 1'd0;
    assign memhint[5519] = 1'd0;
    assign memhint[5520] = 1'd0;
    assign memhint[5521] = 1'd0;
    assign memhint[5522] = 1'd0;
    assign memhint[5523] = 1'd0;
    assign memhint[5524] = 1'd1;
    assign memhint[5525] = 1'd1;
    assign memhint[5526] = 1'd0;
    assign memhint[5527] = 1'd0;
    assign memhint[5528] = 1'd0;
    assign memhint[5529] = 1'd0;
    assign memhint[5530] = 1'd0;
    assign memhint[5531] = 1'd0;
    assign memhint[5532] = 1'd0;
    assign memhint[5533] = 1'd0;
    assign memhint[5534] = 1'd0;
    assign memhint[5535] = 1'd0;
    assign memhint[5536] = 1'd0;
    assign memhint[5537] = 1'd0;
    assign memhint[5538] = 1'd0;
    assign memhint[5539] = 1'd0;
    assign memhint[5540] = 1'd0;
    assign memhint[5541] = 1'd0;
    assign memhint[5542] = 1'd0;
    assign memhint[5543] = 1'd1;
    assign memhint[5544] = 1'd1;
    assign memhint[5545] = 1'd0;
    assign memhint[5546] = 1'd0;
    assign memhint[5547] = 1'd0;
    assign memhint[5548] = 1'd0;
    assign memhint[5549] = 1'd0;
    assign memhint[5550] = 1'd0;
    assign memhint[5551] = 1'd0;
    assign memhint[5552] = 1'd0;
    assign memhint[5553] = 1'd0;
    assign memhint[5554] = 1'd0;
    assign memhint[5555] = 1'd0;
    assign memhint[5556] = 1'd0;
    assign memhint[5557] = 1'd0;
    assign memhint[5558] = 1'd0;
    assign memhint[5559] = 1'd0;
    assign memhint[5560] = 1'd1;
    assign memhint[5561] = 1'd1;
    assign memhint[5562] = 1'd1;
    assign memhint[5563] = 1'd1;
    assign memhint[5564] = 1'd1;
    assign memhint[5565] = 1'd1;
    assign memhint[5566] = 1'd1;
    assign memhint[5567] = 1'd1;
    assign memhint[5568] = 1'd1;
    assign memhint[5569] = 1'd1;
    assign memhint[5570] = 1'd1;
    assign memhint[5571] = 1'd1;
    assign memhint[5572] = 1'd1;
    assign memhint[5573] = 1'd0;
    assign memhint[5574] = 1'd0;
    assign memhint[5575] = 1'd0;
    assign memhint[5576] = 1'd0;
    assign memhint[5577] = 1'd0;
    assign memhint[5578] = 1'd0;
    assign memhint[5579] = 1'd0;
    assign memhint[5580] = 1'd0;
    assign memhint[5581] = 1'd0;
    assign memhint[5582] = 1'd0;
    assign memhint[5583] = 1'd0;
    assign memhint[5584] = 1'd0;
    assign memhint[5585] = 1'd0;
    assign memhint[5586] = 1'd1;
    assign memhint[5587] = 1'd1;
    assign memhint[5588] = 1'd0;
    assign memhint[5589] = 1'd0;
    assign memhint[5590] = 1'd0;
    assign memhint[5591] = 1'd0;
    assign memhint[5592] = 1'd0;
    assign memhint[5593] = 1'd0;
    assign memhint[5594] = 1'd0;
    assign memhint[5595] = 1'd0;
    assign memhint[5596] = 1'd0;
    assign memhint[5597] = 1'd0;
    assign memhint[5598] = 1'd0;
    assign memhint[5599] = 1'd0;
    assign memhint[5600] = 1'd0;
    assign memhint[5601] = 1'd0;
    assign memhint[5602] = 1'd0;
    assign memhint[5603] = 1'd0;
    assign memhint[5604] = 1'd0;
    assign memhint[5605] = 1'd1;
    assign memhint[5606] = 1'd1;
    assign memhint[5607] = 1'd1;
    assign memhint[5608] = 1'd0;
    assign memhint[5609] = 1'd0;
    assign memhint[5610] = 1'd0;
    assign memhint[5611] = 1'd0;
    assign memhint[5612] = 1'd0;
    assign memhint[5613] = 1'd1;
    assign memhint[5614] = 1'd1;
    assign memhint[5615] = 1'd0;
    assign memhint[5616] = 1'd0;
    assign memhint[5617] = 1'd0;
    assign memhint[5618] = 1'd0;
    assign memhint[5619] = 1'd0;
    assign memhint[5620] = 1'd0;
    assign memhint[5621] = 1'd0;
    assign memhint[5622] = 1'd0;
    assign memhint[5623] = 1'd0;
    assign memhint[5624] = 1'd0;
    assign memhint[5625] = 1'd0;
    assign memhint[5626] = 1'd0;
    assign memhint[5627] = 1'd0;
    assign memhint[5628] = 1'd0;
    assign memhint[5629] = 1'd0;
    assign memhint[5630] = 1'd1;
    assign memhint[5631] = 1'd1;
    assign memhint[5632] = 1'd0;
    assign memhint[5633] = 1'd0;
    assign memhint[5634] = 1'd0;
    assign memhint[5635] = 1'd0;
    assign memhint[5636] = 1'd0;
    assign memhint[5637] = 1'd0;
    assign memhint[5638] = 1'd0;
    assign memhint[5639] = 1'd0;
    assign memhint[5640] = 1'd0;
    assign memhint[5641] = 1'd0;
    assign memhint[5642] = 1'd0;
    assign memhint[5643] = 1'd0;
    assign memhint[5644] = 1'd0;
    assign memhint[5645] = 1'd1;
    assign memhint[5646] = 1'd1;
    assign memhint[5647] = 1'd0;
    assign memhint[5648] = 1'd0;
    assign memhint[5649] = 1'd0;
    assign memhint[5650] = 1'd0;
    assign memhint[5651] = 1'd0;
    assign memhint[5652] = 1'd0;
    assign memhint[5653] = 1'd0;
    assign memhint[5654] = 1'd0;
    assign memhint[5655] = 1'd0;
    assign memhint[5656] = 1'd0;
    assign memhint[5657] = 1'd0;
    assign memhint[5658] = 1'd0;
    assign memhint[5659] = 1'd0;
    assign memhint[5660] = 1'd0;
    assign memhint[5661] = 1'd0;
    assign memhint[5662] = 1'd1;
    assign memhint[5663] = 1'd1;
    assign memhint[5664] = 1'd0;
    assign memhint[5665] = 1'd0;
    assign memhint[5666] = 1'd0;
    assign memhint[5667] = 1'd0;
    assign memhint[5668] = 1'd0;
    assign memhint[5669] = 1'd0;
    assign memhint[5670] = 1'd0;
    assign memhint[5671] = 1'd0;
    assign memhint[5672] = 1'd0;
    assign memhint[5673] = 1'd0;
    assign memhint[5674] = 1'd0;
    assign memhint[5675] = 1'd0;
    assign memhint[5676] = 1'd0;
    assign memhint[5677] = 1'd0;
    assign memhint[5678] = 1'd0;
    assign memhint[5679] = 1'd0;
    assign memhint[5680] = 1'd0;
    assign memhint[5681] = 1'd0;
    assign memhint[5682] = 1'd0;
    assign memhint[5683] = 1'd0;
    assign memhint[5684] = 1'd0;
    assign memhint[5685] = 1'd0;
    assign memhint[5686] = 1'd0;
    assign memhint[5687] = 1'd0;
    assign memhint[5688] = 1'd0;
    assign memhint[5689] = 1'd0;
    assign memhint[5690] = 1'd1;
    assign memhint[5691] = 1'd1;
    assign memhint[5692] = 1'd0;
    assign memhint[5693] = 1'd0;
    assign memhint[5694] = 1'd0;
    assign memhint[5695] = 1'd0;
    assign memhint[5696] = 1'd0;
    assign memhint[5697] = 1'd0;
    assign memhint[5698] = 1'd0;
    assign memhint[5699] = 1'd0;
    assign memhint[5700] = 1'd0;
    assign memhint[5701] = 1'd0;
    assign memhint[5702] = 1'd0;
    assign memhint[5703] = 1'd0;
    assign memhint[5704] = 1'd0;
    assign memhint[5705] = 1'd0;
    assign memhint[5706] = 1'd0;
    assign memhint[5707] = 1'd0;
    assign memhint[5708] = 1'd0;
    assign memhint[5709] = 1'd0;
    assign memhint[5710] = 1'd0;
    assign memhint[5711] = 1'd1;
    assign memhint[5712] = 1'd1;
    assign memhint[5713] = 1'd0;
    assign memhint[5714] = 1'd0;
    assign memhint[5715] = 1'd0;
    assign memhint[5716] = 1'd0;
    assign memhint[5717] = 1'd0;
    assign memhint[5718] = 1'd0;
    assign memhint[5719] = 1'd0;
    assign memhint[5720] = 1'd0;
    assign memhint[5721] = 1'd0;
    assign memhint[5722] = 1'd0;
    assign memhint[5723] = 1'd0;
    assign memhint[5724] = 1'd1;
    assign memhint[5725] = 1'd1;
    assign memhint[5726] = 1'd0;
    assign memhint[5727] = 1'd0;
    assign memhint[5728] = 1'd0;
    assign memhint[5729] = 1'd0;
    assign memhint[5730] = 1'd0;
    assign memhint[5731] = 1'd0;
    assign memhint[5732] = 1'd0;
    assign memhint[5733] = 1'd0;
    assign memhint[5734] = 1'd0;
    assign memhint[5735] = 1'd0;
    assign memhint[5736] = 1'd0;
    assign memhint[5737] = 1'd0;
    assign memhint[5738] = 1'd0;
    assign memhint[5739] = 1'd0;
    assign memhint[5740] = 1'd0;
    assign memhint[5741] = 1'd0;
    assign memhint[5742] = 1'd0;
    assign memhint[5743] = 1'd0;
    assign memhint[5744] = 1'd0;
    assign memhint[5745] = 1'd0;
    assign memhint[5746] = 1'd0;
    assign memhint[5747] = 1'd0;
    assign memhint[5748] = 1'd0;
    assign memhint[5749] = 1'd0;
    assign memhint[5750] = 1'd1;
    assign memhint[5751] = 1'd1;
    assign memhint[5752] = 1'd1;
    assign memhint[5753] = 1'd0;
    assign memhint[5754] = 1'd0;
    assign memhint[5755] = 1'd0;
    assign memhint[5756] = 1'd0;
    assign memhint[5757] = 1'd0;
    assign memhint[5758] = 1'd1;
    assign memhint[5759] = 1'd1;
    assign memhint[5760] = 1'd0;
    assign memhint[5761] = 1'd0;
    assign memhint[5762] = 1'd0;
    assign memhint[5763] = 1'd0;
    assign memhint[5764] = 1'd0;
    assign memhint[5765] = 1'd0;
    assign memhint[5766] = 1'd0;
    assign memhint[5767] = 1'd0;
    assign memhint[5768] = 1'd0;
    assign memhint[5769] = 1'd0;
    assign memhint[5770] = 1'd0;
    assign memhint[5771] = 1'd0;
    assign memhint[5772] = 1'd0;
    assign memhint[5773] = 1'd0;
    assign memhint[5774] = 1'd0;
    assign memhint[5775] = 1'd0;
    assign memhint[5776] = 1'd0;
    assign memhint[5777] = 1'd0;
    assign memhint[5778] = 1'd1;
    assign memhint[5779] = 1'd1;
    assign memhint[5780] = 1'd0;
    assign memhint[5781] = 1'd0;
    assign memhint[5782] = 1'd0;
    assign memhint[5783] = 1'd0;
    assign memhint[5784] = 1'd0;
    assign memhint[5785] = 1'd0;
    assign memhint[5786] = 1'd1;
    assign memhint[5787] = 1'd1;
    assign memhint[5788] = 1'd0;
    assign memhint[5789] = 1'd0;
    assign memhint[5790] = 1'd0;
    assign memhint[5791] = 1'd0;
    assign memhint[5792] = 1'd0;
    assign memhint[5793] = 1'd0;
    assign memhint[5794] = 1'd0;
    assign memhint[5795] = 1'd0;
    assign memhint[5796] = 1'd0;
    assign memhint[5797] = 1'd1;
    assign memhint[5798] = 1'd1;
    assign memhint[5799] = 1'd0;
    assign memhint[5800] = 1'd0;
    assign memhint[5801] = 1'd0;
    assign memhint[5802] = 1'd1;
    assign memhint[5803] = 1'd1;
    assign memhint[5804] = 1'd0;
    assign memhint[5805] = 1'd0;
    assign memhint[5806] = 1'd0;
    assign memhint[5807] = 1'd0;
    assign memhint[5808] = 1'd0;
    assign memhint[5809] = 1'd0;
    assign memhint[5810] = 1'd1;
    assign memhint[5811] = 1'd1;
    assign memhint[5812] = 1'd0;
    assign memhint[5813] = 1'd0;
    assign memhint[5814] = 1'd0;
    assign memhint[5815] = 1'd0;
    assign memhint[5816] = 1'd0;
    assign memhint[5817] = 1'd0;
    assign memhint[5818] = 1'd0;
    assign memhint[5819] = 1'd0;
    assign memhint[5820] = 1'd0;
    assign memhint[5821] = 1'd0;
    assign memhint[5822] = 1'd0;
    assign memhint[5823] = 1'd0;
    assign memhint[5824] = 1'd0;
    assign memhint[5825] = 1'd0;
    assign memhint[5826] = 1'd0;
    assign memhint[5827] = 1'd0;
    assign memhint[5828] = 1'd0;
    assign memhint[5829] = 1'd0;
    assign memhint[5830] = 1'd0;
    assign memhint[5831] = 1'd1;
    assign memhint[5832] = 1'd1;
    assign memhint[5833] = 1'd0;
    assign memhint[5834] = 1'd0;
    assign memhint[5835] = 1'd0;
    assign memhint[5836] = 1'd0;
    assign memhint[5837] = 1'd0;
    assign memhint[5838] = 1'd0;
    assign memhint[5839] = 1'd0;
    assign memhint[5840] = 1'd0;
    assign memhint[5841] = 1'd0;
    assign memhint[5842] = 1'd0;
    assign memhint[5843] = 1'd0;
    assign memhint[5844] = 1'd0;
    assign memhint[5845] = 1'd0;
    assign memhint[5846] = 1'd0;
    assign memhint[5847] = 1'd0;
    assign memhint[5848] = 1'd0;
    assign memhint[5849] = 1'd1;
    assign memhint[5850] = 1'd1;
    assign memhint[5851] = 1'd0;
    assign memhint[5852] = 1'd0;
    assign memhint[5853] = 1'd0;
    assign memhint[5854] = 1'd0;
    assign memhint[5855] = 1'd0;
    assign memhint[5856] = 1'd0;
    assign memhint[5857] = 1'd0;
    assign memhint[5858] = 1'd0;
    assign memhint[5859] = 1'd0;
    assign memhint[5860] = 1'd1;
    assign memhint[5861] = 1'd1;
    assign memhint[5862] = 1'd0;
    assign memhint[5863] = 1'd0;
    assign memhint[5864] = 1'd0;
    assign memhint[5865] = 1'd0;
    assign memhint[5866] = 1'd0;
    assign memhint[5867] = 1'd0;
    assign memhint[5868] = 1'd0;
    assign memhint[5869] = 1'd0;
    assign memhint[5870] = 1'd0;
    assign memhint[5871] = 1'd0;
    assign memhint[5872] = 1'd0;
    assign memhint[5873] = 1'd0;
    assign memhint[5874] = 1'd0;
    assign memhint[5875] = 1'd0;
    assign memhint[5876] = 1'd0;
    assign memhint[5877] = 1'd0;
    assign memhint[5878] = 1'd0;
    assign memhint[5879] = 1'd0;
    assign memhint[5880] = 1'd1;
    assign memhint[5881] = 1'd1;
    assign memhint[5882] = 1'd0;
    assign memhint[5883] = 1'd0;
    assign memhint[5884] = 1'd0;
    assign memhint[5885] = 1'd0;
    assign memhint[5886] = 1'd0;
    assign memhint[5887] = 1'd0;
    assign memhint[5888] = 1'd0;
    assign memhint[5889] = 1'd0;
    assign memhint[5890] = 1'd0;
    assign memhint[5891] = 1'd0;
    assign memhint[5892] = 1'd0;
    assign memhint[5893] = 1'd0;
    assign memhint[5894] = 1'd0;
    assign memhint[5895] = 1'd0;
    assign memhint[5896] = 1'd0;
    assign memhint[5897] = 1'd1;
    assign memhint[5898] = 1'd1;
    assign memhint[5899] = 1'd0;
    assign memhint[5900] = 1'd0;
    assign memhint[5901] = 1'd0;
    assign memhint[5902] = 1'd0;
    assign memhint[5903] = 1'd0;
    assign memhint[5904] = 1'd0;
    assign memhint[5905] = 1'd0;
    assign memhint[5906] = 1'd0;
    assign memhint[5907] = 1'd0;
    assign memhint[5908] = 1'd0;
    assign memhint[5909] = 1'd0;
    assign memhint[5910] = 1'd0;
    assign memhint[5911] = 1'd0;
    assign memhint[5912] = 1'd0;
    assign memhint[5913] = 1'd0;
    assign memhint[5914] = 1'd0;
    assign memhint[5915] = 1'd0;
    assign memhint[5916] = 1'd1;
    assign memhint[5917] = 1'd1;
    assign memhint[5918] = 1'd0;
    assign memhint[5919] = 1'd0;
    assign memhint[5920] = 1'd0;
    assign memhint[5921] = 1'd0;
    assign memhint[5922] = 1'd0;
    assign memhint[5923] = 1'd0;
    assign memhint[5924] = 1'd0;
    assign memhint[5925] = 1'd0;
    assign memhint[5926] = 1'd0;
    assign memhint[5927] = 1'd0;
    assign memhint[5928] = 1'd0;
    assign memhint[5929] = 1'd0;
    assign memhint[5930] = 1'd0;
    assign memhint[5931] = 1'd0;
    assign memhint[5932] = 1'd1;
    assign memhint[5933] = 1'd1;
    assign memhint[5934] = 1'd0;
    assign memhint[5935] = 1'd0;
    assign memhint[5936] = 1'd0;
    assign memhint[5937] = 1'd0;
    assign memhint[5938] = 1'd0;
    assign memhint[5939] = 1'd0;
    assign memhint[5940] = 1'd0;
    assign memhint[5941] = 1'd0;
    assign memhint[5942] = 1'd0;
    assign memhint[5943] = 1'd0;
    assign memhint[5944] = 1'd0;
    assign memhint[5945] = 1'd1;
    assign memhint[5946] = 1'd1;
    assign memhint[5947] = 1'd0;
    assign memhint[5948] = 1'd0;
    assign memhint[5949] = 1'd0;
    assign memhint[5950] = 1'd0;
    assign memhint[5951] = 1'd0;
    assign memhint[5952] = 1'd0;
    assign memhint[5953] = 1'd0;
    assign memhint[5954] = 1'd0;
    assign memhint[5955] = 1'd0;
    assign memhint[5956] = 1'd0;
    assign memhint[5957] = 1'd0;
    assign memhint[5958] = 1'd0;
    assign memhint[5959] = 1'd1;
    assign memhint[5960] = 1'd1;
    assign memhint[5961] = 1'd0;
    assign memhint[5962] = 1'd0;
    assign memhint[5963] = 1'd0;
    assign memhint[5964] = 1'd0;
    assign memhint[5965] = 1'd0;
    assign memhint[5966] = 1'd0;
    assign memhint[5967] = 1'd0;
    assign memhint[5968] = 1'd0;
    assign memhint[5969] = 1'd0;
    assign memhint[5970] = 1'd0;
    assign memhint[5971] = 1'd0;
    assign memhint[5972] = 1'd0;
    assign memhint[5973] = 1'd0;
    assign memhint[5974] = 1'd0;
    assign memhint[5975] = 1'd0;
    assign memhint[5976] = 1'd0;
    assign memhint[5977] = 1'd0;
    assign memhint[5978] = 1'd0;
    assign memhint[5979] = 1'd1;
    assign memhint[5980] = 1'd1;
    assign memhint[5981] = 1'd0;
    assign memhint[5982] = 1'd0;
    assign memhint[5983] = 1'd0;
    assign memhint[5984] = 1'd0;
    assign memhint[5985] = 1'd0;
    assign memhint[5986] = 1'd1;
    assign memhint[5987] = 1'd1;
    assign memhint[5988] = 1'd0;
    assign memhint[5989] = 1'd0;
    assign memhint[5990] = 1'd0;
    assign memhint[5991] = 1'd0;
    assign memhint[5992] = 1'd0;
    assign memhint[5993] = 1'd0;
    assign memhint[5994] = 1'd0;
    assign memhint[5995] = 1'd0;
    assign memhint[5996] = 1'd0;
    assign memhint[5997] = 1'd0;
    assign memhint[5998] = 1'd0;
    assign memhint[5999] = 1'd0;
    assign memhint[6000] = 1'd0;
    assign memhint[6001] = 1'd0;
    assign memhint[6002] = 1'd0;
    assign memhint[6003] = 1'd1;
    assign memhint[6004] = 1'd1;
    assign memhint[6005] = 1'd0;
    assign memhint[6006] = 1'd0;
    assign memhint[6007] = 1'd0;
    assign memhint[6008] = 1'd0;
    assign memhint[6009] = 1'd0;
    assign memhint[6010] = 1'd0;
    assign memhint[6011] = 1'd0;
    assign memhint[6012] = 1'd0;
    assign memhint[6013] = 1'd0;
    assign memhint[6014] = 1'd0;
    assign memhint[6015] = 1'd0;
    assign memhint[6016] = 1'd0;
    assign memhint[6017] = 1'd0;
    assign memhint[6018] = 1'd1;
    assign memhint[6019] = 1'd1;
    assign memhint[6020] = 1'd0;
    assign memhint[6021] = 1'd0;
    assign memhint[6022] = 1'd0;
    assign memhint[6023] = 1'd0;
    assign memhint[6024] = 1'd0;
    assign memhint[6025] = 1'd0;
    assign memhint[6026] = 1'd0;
    assign memhint[6027] = 1'd0;
    assign memhint[6028] = 1'd0;
    assign memhint[6029] = 1'd0;
    assign memhint[6030] = 1'd0;
    assign memhint[6031] = 1'd0;
    assign memhint[6032] = 1'd0;
    assign memhint[6033] = 1'd0;
    assign memhint[6034] = 1'd0;
    assign memhint[6035] = 1'd1;
    assign memhint[6036] = 1'd1;
    assign memhint[6037] = 1'd0;
    assign memhint[6038] = 1'd0;
    assign memhint[6039] = 1'd0;
    assign memhint[6040] = 1'd0;
    assign memhint[6041] = 1'd0;
    assign memhint[6042] = 1'd0;
    assign memhint[6043] = 1'd0;
    assign memhint[6044] = 1'd0;
    assign memhint[6045] = 1'd0;
    assign memhint[6046] = 1'd0;
    assign memhint[6047] = 1'd0;
    assign memhint[6048] = 1'd0;
    assign memhint[6049] = 1'd0;
    assign memhint[6050] = 1'd0;
    assign memhint[6051] = 1'd0;
    assign memhint[6052] = 1'd0;
    assign memhint[6053] = 1'd0;
    assign memhint[6054] = 1'd0;
    assign memhint[6055] = 1'd0;
    assign memhint[6056] = 1'd0;
    assign memhint[6057] = 1'd0;
    assign memhint[6058] = 1'd0;
    assign memhint[6059] = 1'd0;
    assign memhint[6060] = 1'd0;
    assign memhint[6061] = 1'd0;
    assign memhint[6062] = 1'd0;
    assign memhint[6063] = 1'd1;
    assign memhint[6064] = 1'd1;
    assign memhint[6065] = 1'd0;
    assign memhint[6066] = 1'd0;
    assign memhint[6067] = 1'd0;
    assign memhint[6068] = 1'd0;
    assign memhint[6069] = 1'd0;
    assign memhint[6070] = 1'd0;
    assign memhint[6071] = 1'd0;
    assign memhint[6072] = 1'd0;
    assign memhint[6073] = 1'd0;
    assign memhint[6074] = 1'd0;
    assign memhint[6075] = 1'd0;
    assign memhint[6076] = 1'd0;
    assign memhint[6077] = 1'd0;
    assign memhint[6078] = 1'd0;
    assign memhint[6079] = 1'd0;
    assign memhint[6080] = 1'd0;
    assign memhint[6081] = 1'd0;
    assign memhint[6082] = 1'd0;
    assign memhint[6083] = 1'd0;
    assign memhint[6084] = 1'd1;
    assign memhint[6085] = 1'd1;
    assign memhint[6086] = 1'd0;
    assign memhint[6087] = 1'd0;
    assign memhint[6088] = 1'd0;
    assign memhint[6089] = 1'd0;
    assign memhint[6090] = 1'd0;
    assign memhint[6091] = 1'd0;
    assign memhint[6092] = 1'd0;
    assign memhint[6093] = 1'd0;
    assign memhint[6094] = 1'd0;
    assign memhint[6095] = 1'd0;
    assign memhint[6096] = 1'd0;
    assign memhint[6097] = 1'd1;
    assign memhint[6098] = 1'd1;
    assign memhint[6099] = 1'd0;
    assign memhint[6100] = 1'd0;
    assign memhint[6101] = 1'd0;
    assign memhint[6102] = 1'd0;
    assign memhint[6103] = 1'd0;
    assign memhint[6104] = 1'd0;
    assign memhint[6105] = 1'd0;
    assign memhint[6106] = 1'd0;
    assign memhint[6107] = 1'd0;
    assign memhint[6108] = 1'd0;
    assign memhint[6109] = 1'd0;
    assign memhint[6110] = 1'd0;
    assign memhint[6111] = 1'd0;
    assign memhint[6112] = 1'd0;
    assign memhint[6113] = 1'd0;
    assign memhint[6114] = 1'd0;
    assign memhint[6115] = 1'd0;
    assign memhint[6116] = 1'd0;
    assign memhint[6117] = 1'd0;
    assign memhint[6118] = 1'd0;
    assign memhint[6119] = 1'd0;
    assign memhint[6120] = 1'd0;
    assign memhint[6121] = 1'd0;
    assign memhint[6122] = 1'd0;
    assign memhint[6123] = 1'd0;
    assign memhint[6124] = 1'd1;
    assign memhint[6125] = 1'd1;
    assign memhint[6126] = 1'd0;
    assign memhint[6127] = 1'd0;
    assign memhint[6128] = 1'd0;
    assign memhint[6129] = 1'd0;
    assign memhint[6130] = 1'd0;
    assign memhint[6131] = 1'd1;
    assign memhint[6132] = 1'd1;
    assign memhint[6133] = 1'd0;
    assign memhint[6134] = 1'd0;
    assign memhint[6135] = 1'd0;
    assign memhint[6136] = 1'd0;
    assign memhint[6137] = 1'd0;
    assign memhint[6138] = 1'd0;
    assign memhint[6139] = 1'd0;
    assign memhint[6140] = 1'd0;
    assign memhint[6141] = 1'd0;
    assign memhint[6142] = 1'd0;
    assign memhint[6143] = 1'd0;
    assign memhint[6144] = 1'd0;
    assign memhint[6145] = 1'd0;
    assign memhint[6146] = 1'd0;
    assign memhint[6147] = 1'd0;
    assign memhint[6148] = 1'd0;
    assign memhint[6149] = 1'd0;
    assign memhint[6150] = 1'd0;
    assign memhint[6151] = 1'd1;
    assign memhint[6152] = 1'd1;
    assign memhint[6153] = 1'd0;
    assign memhint[6154] = 1'd0;
    assign memhint[6155] = 1'd0;
    assign memhint[6156] = 1'd0;
    assign memhint[6157] = 1'd0;
    assign memhint[6158] = 1'd0;
    assign memhint[6159] = 1'd1;
    assign memhint[6160] = 1'd1;
    assign memhint[6161] = 1'd0;
    assign memhint[6162] = 1'd0;
    assign memhint[6163] = 1'd0;
    assign memhint[6164] = 1'd0;
    assign memhint[6165] = 1'd0;
    assign memhint[6166] = 1'd0;
    assign memhint[6167] = 1'd0;
    assign memhint[6168] = 1'd0;
    assign memhint[6169] = 1'd0;
    assign memhint[6170] = 1'd0;
    assign memhint[6171] = 1'd1;
    assign memhint[6172] = 1'd1;
    assign memhint[6173] = 1'd0;
    assign memhint[6174] = 1'd0;
    assign memhint[6175] = 1'd1;
    assign memhint[6176] = 1'd1;
    assign memhint[6177] = 1'd0;
    assign memhint[6178] = 1'd0;
    assign memhint[6179] = 1'd0;
    assign memhint[6180] = 1'd0;
    assign memhint[6181] = 1'd0;
    assign memhint[6182] = 1'd0;
    assign memhint[6183] = 1'd1;
    assign memhint[6184] = 1'd1;
    assign memhint[6185] = 1'd1;
    assign memhint[6186] = 1'd0;
    assign memhint[6187] = 1'd0;
    assign memhint[6188] = 1'd0;
    assign memhint[6189] = 1'd0;
    assign memhint[6190] = 1'd0;
    assign memhint[6191] = 1'd0;
    assign memhint[6192] = 1'd0;
    assign memhint[6193] = 1'd0;
    assign memhint[6194] = 1'd0;
    assign memhint[6195] = 1'd0;
    assign memhint[6196] = 1'd0;
    assign memhint[6197] = 1'd0;
    assign memhint[6198] = 1'd0;
    assign memhint[6199] = 1'd0;
    assign memhint[6200] = 1'd0;
    assign memhint[6201] = 1'd0;
    assign memhint[6202] = 1'd0;
    assign memhint[6203] = 1'd1;
    assign memhint[6204] = 1'd1;
    assign memhint[6205] = 1'd0;
    assign memhint[6206] = 1'd0;
    assign memhint[6207] = 1'd0;
    assign memhint[6208] = 1'd0;
    assign memhint[6209] = 1'd0;
    assign memhint[6210] = 1'd0;
    assign memhint[6211] = 1'd0;
    assign memhint[6212] = 1'd0;
    assign memhint[6213] = 1'd0;
    assign memhint[6214] = 1'd0;
    assign memhint[6215] = 1'd0;
    assign memhint[6216] = 1'd0;
    assign memhint[6217] = 1'd0;
    assign memhint[6218] = 1'd0;
    assign memhint[6219] = 1'd0;
    assign memhint[6220] = 1'd0;
    assign memhint[6221] = 1'd0;
    assign memhint[6222] = 1'd1;
    assign memhint[6223] = 1'd1;
    assign memhint[6224] = 1'd0;
    assign memhint[6225] = 1'd0;
    assign memhint[6226] = 1'd0;
    assign memhint[6227] = 1'd0;
    assign memhint[6228] = 1'd0;
    assign memhint[6229] = 1'd0;
    assign memhint[6230] = 1'd0;
    assign memhint[6231] = 1'd0;
    assign memhint[6232] = 1'd0;
    assign memhint[6233] = 1'd1;
    assign memhint[6234] = 1'd1;
    assign memhint[6235] = 1'd0;
    assign memhint[6236] = 1'd0;
    assign memhint[6237] = 1'd0;
    assign memhint[6238] = 1'd0;
    assign memhint[6239] = 1'd0;
    assign memhint[6240] = 1'd0;
    assign memhint[6241] = 1'd0;
    assign memhint[6242] = 1'd0;
    assign memhint[6243] = 1'd0;
    assign memhint[6244] = 1'd0;
    assign memhint[6245] = 1'd0;
    assign memhint[6246] = 1'd0;
    assign memhint[6247] = 1'd0;
    assign memhint[6248] = 1'd0;
    assign memhint[6249] = 1'd0;
    assign memhint[6250] = 1'd0;
    assign memhint[6251] = 1'd0;
    assign memhint[6252] = 1'd0;
    assign memhint[6253] = 1'd1;
    assign memhint[6254] = 1'd1;
    assign memhint[6255] = 1'd0;
    assign memhint[6256] = 1'd0;
    assign memhint[6257] = 1'd0;
    assign memhint[6258] = 1'd0;
    assign memhint[6259] = 1'd0;
    assign memhint[6260] = 1'd0;
    assign memhint[6261] = 1'd0;
    assign memhint[6262] = 1'd0;
    assign memhint[6263] = 1'd0;
    assign memhint[6264] = 1'd0;
    assign memhint[6265] = 1'd0;
    assign memhint[6266] = 1'd0;
    assign memhint[6267] = 1'd0;
    assign memhint[6268] = 1'd0;
    assign memhint[6269] = 1'd0;
    assign memhint[6270] = 1'd1;
    assign memhint[6271] = 1'd1;
    assign memhint[6272] = 1'd0;
    assign memhint[6273] = 1'd0;
    assign memhint[6274] = 1'd0;
    assign memhint[6275] = 1'd0;
    assign memhint[6276] = 1'd0;
    assign memhint[6277] = 1'd0;
    assign memhint[6278] = 1'd0;
    assign memhint[6279] = 1'd0;
    assign memhint[6280] = 1'd0;
    assign memhint[6281] = 1'd0;
    assign memhint[6282] = 1'd0;
    assign memhint[6283] = 1'd0;
    assign memhint[6284] = 1'd0;
    assign memhint[6285] = 1'd0;
    assign memhint[6286] = 1'd0;
    assign memhint[6287] = 1'd0;
    assign memhint[6288] = 1'd0;
    assign memhint[6289] = 1'd1;
    assign memhint[6290] = 1'd1;
    assign memhint[6291] = 1'd0;
    assign memhint[6292] = 1'd0;
    assign memhint[6293] = 1'd0;
    assign memhint[6294] = 1'd0;
    assign memhint[6295] = 1'd0;
    assign memhint[6296] = 1'd0;
    assign memhint[6297] = 1'd0;
    assign memhint[6298] = 1'd0;
    assign memhint[6299] = 1'd0;
    assign memhint[6300] = 1'd0;
    assign memhint[6301] = 1'd0;
    assign memhint[6302] = 1'd0;
    assign memhint[6303] = 1'd0;
    assign memhint[6304] = 1'd0;
    assign memhint[6305] = 1'd1;
    assign memhint[6306] = 1'd1;
    assign memhint[6307] = 1'd0;
    assign memhint[6308] = 1'd0;
    assign memhint[6309] = 1'd0;
    assign memhint[6310] = 1'd0;
    assign memhint[6311] = 1'd0;
    assign memhint[6312] = 1'd0;
    assign memhint[6313] = 1'd0;
    assign memhint[6314] = 1'd0;
    assign memhint[6315] = 1'd0;
    assign memhint[6316] = 1'd0;
    assign memhint[6317] = 1'd0;
    assign memhint[6318] = 1'd1;
    assign memhint[6319] = 1'd1;
    assign memhint[6320] = 1'd0;
    assign memhint[6321] = 1'd0;
    assign memhint[6322] = 1'd0;
    assign memhint[6323] = 1'd0;
    assign memhint[6324] = 1'd0;
    assign memhint[6325] = 1'd0;
    assign memhint[6326] = 1'd0;
    assign memhint[6327] = 1'd0;
    assign memhint[6328] = 1'd0;
    assign memhint[6329] = 1'd0;
    assign memhint[6330] = 1'd0;
    assign memhint[6331] = 1'd0;
    assign memhint[6332] = 1'd1;
    assign memhint[6333] = 1'd1;
    assign memhint[6334] = 1'd0;
    assign memhint[6335] = 1'd0;
    assign memhint[6336] = 1'd0;
    assign memhint[6337] = 1'd0;
    assign memhint[6338] = 1'd0;
    assign memhint[6339] = 1'd0;
    assign memhint[6340] = 1'd0;
    assign memhint[6341] = 1'd0;
    assign memhint[6342] = 1'd1;
    assign memhint[6343] = 1'd0;
    assign memhint[6344] = 1'd0;
    assign memhint[6345] = 1'd0;
    assign memhint[6346] = 1'd0;
    assign memhint[6347] = 1'd0;
    assign memhint[6348] = 1'd0;
    assign memhint[6349] = 1'd0;
    assign memhint[6350] = 1'd0;
    assign memhint[6351] = 1'd0;
    assign memhint[6352] = 1'd1;
    assign memhint[6353] = 1'd1;
    assign memhint[6354] = 1'd0;
    assign memhint[6355] = 1'd0;
    assign memhint[6356] = 1'd0;
    assign memhint[6357] = 1'd0;
    assign memhint[6358] = 1'd0;
    assign memhint[6359] = 1'd1;
    assign memhint[6360] = 1'd1;
    assign memhint[6361] = 1'd0;
    assign memhint[6362] = 1'd0;
    assign memhint[6363] = 1'd0;
    assign memhint[6364] = 1'd0;
    assign memhint[6365] = 1'd0;
    assign memhint[6366] = 1'd0;
    assign memhint[6367] = 1'd0;
    assign memhint[6368] = 1'd0;
    assign memhint[6369] = 1'd0;
    assign memhint[6370] = 1'd0;
    assign memhint[6371] = 1'd0;
    assign memhint[6372] = 1'd0;
    assign memhint[6373] = 1'd0;
    assign memhint[6374] = 1'd0;
    assign memhint[6375] = 1'd0;
    assign memhint[6376] = 1'd1;
    assign memhint[6377] = 1'd1;
    assign memhint[6378] = 1'd0;
    assign memhint[6379] = 1'd0;
    assign memhint[6380] = 1'd0;
    assign memhint[6381] = 1'd0;
    assign memhint[6382] = 1'd0;
    assign memhint[6383] = 1'd0;
    assign memhint[6384] = 1'd0;
    assign memhint[6385] = 1'd0;
    assign memhint[6386] = 1'd0;
    assign memhint[6387] = 1'd0;
    assign memhint[6388] = 1'd0;
    assign memhint[6389] = 1'd0;
    assign memhint[6390] = 1'd0;
    assign memhint[6391] = 1'd1;
    assign memhint[6392] = 1'd1;
    assign memhint[6393] = 1'd0;
    assign memhint[6394] = 1'd0;
    assign memhint[6395] = 1'd0;
    assign memhint[6396] = 1'd0;
    assign memhint[6397] = 1'd0;
    assign memhint[6398] = 1'd0;
    assign memhint[6399] = 1'd0;
    assign memhint[6400] = 1'd0;
    assign memhint[6401] = 1'd0;
    assign memhint[6402] = 1'd0;
    assign memhint[6403] = 1'd0;
    assign memhint[6404] = 1'd0;
    assign memhint[6405] = 1'd0;
    assign memhint[6406] = 1'd0;
    assign memhint[6407] = 1'd0;
    assign memhint[6408] = 1'd0;
    assign memhint[6409] = 1'd1;
    assign memhint[6410] = 1'd1;
    assign memhint[6411] = 1'd0;
    assign memhint[6412] = 1'd0;
    assign memhint[6413] = 1'd0;
    assign memhint[6414] = 1'd0;
    assign memhint[6415] = 1'd0;
    assign memhint[6416] = 1'd0;
    assign memhint[6417] = 1'd0;
    assign memhint[6418] = 1'd0;
    assign memhint[6419] = 1'd0;
    assign memhint[6420] = 1'd0;
    assign memhint[6421] = 1'd0;
    assign memhint[6422] = 1'd0;
    assign memhint[6423] = 1'd0;
    assign memhint[6424] = 1'd0;
    assign memhint[6425] = 1'd0;
    assign memhint[6426] = 1'd0;
    assign memhint[6427] = 1'd1;
    assign memhint[6428] = 1'd0;
    assign memhint[6429] = 1'd0;
    assign memhint[6430] = 1'd0;
    assign memhint[6431] = 1'd0;
    assign memhint[6432] = 1'd0;
    assign memhint[6433] = 1'd0;
    assign memhint[6434] = 1'd0;
    assign memhint[6435] = 1'd0;
    assign memhint[6436] = 1'd1;
    assign memhint[6437] = 1'd1;
    assign memhint[6438] = 1'd0;
    assign memhint[6439] = 1'd0;
    assign memhint[6440] = 1'd0;
    assign memhint[6441] = 1'd0;
    assign memhint[6442] = 1'd0;
    assign memhint[6443] = 1'd0;
    assign memhint[6444] = 1'd0;
    assign memhint[6445] = 1'd0;
    assign memhint[6446] = 1'd0;
    assign memhint[6447] = 1'd0;
    assign memhint[6448] = 1'd0;
    assign memhint[6449] = 1'd0;
    assign memhint[6450] = 1'd0;
    assign memhint[6451] = 1'd0;
    assign memhint[6452] = 1'd0;
    assign memhint[6453] = 1'd0;
    assign memhint[6454] = 1'd0;
    assign memhint[6455] = 1'd0;
    assign memhint[6456] = 1'd1;
    assign memhint[6457] = 1'd1;
    assign memhint[6458] = 1'd1;
    assign memhint[6459] = 1'd0;
    assign memhint[6460] = 1'd0;
    assign memhint[6461] = 1'd0;
    assign memhint[6462] = 1'd0;
    assign memhint[6463] = 1'd0;
    assign memhint[6464] = 1'd0;
    assign memhint[6465] = 1'd0;
    assign memhint[6466] = 1'd0;
    assign memhint[6467] = 1'd0;
    assign memhint[6468] = 1'd0;
    assign memhint[6469] = 1'd0;
    assign memhint[6470] = 1'd0;
    assign memhint[6471] = 1'd1;
    assign memhint[6472] = 1'd1;
    assign memhint[6473] = 1'd0;
    assign memhint[6474] = 1'd0;
    assign memhint[6475] = 1'd0;
    assign memhint[6476] = 1'd0;
    assign memhint[6477] = 1'd0;
    assign memhint[6478] = 1'd0;
    assign memhint[6479] = 1'd0;
    assign memhint[6480] = 1'd0;
    assign memhint[6481] = 1'd0;
    assign memhint[6482] = 1'd0;
    assign memhint[6483] = 1'd0;
    assign memhint[6484] = 1'd0;
    assign memhint[6485] = 1'd0;
    assign memhint[6486] = 1'd0;
    assign memhint[6487] = 1'd1;
    assign memhint[6488] = 1'd0;
    assign memhint[6489] = 1'd0;
    assign memhint[6490] = 1'd0;
    assign memhint[6491] = 1'd0;
    assign memhint[6492] = 1'd0;
    assign memhint[6493] = 1'd0;
    assign memhint[6494] = 1'd0;
    assign memhint[6495] = 1'd0;
    assign memhint[6496] = 1'd0;
    assign memhint[6497] = 1'd1;
    assign memhint[6498] = 1'd1;
    assign memhint[6499] = 1'd0;
    assign memhint[6500] = 1'd0;
    assign memhint[6501] = 1'd0;
    assign memhint[6502] = 1'd0;
    assign memhint[6503] = 1'd0;
    assign memhint[6504] = 1'd0;
    assign memhint[6505] = 1'd1;
    assign memhint[6506] = 1'd1;
    assign memhint[6507] = 1'd0;
    assign memhint[6508] = 1'd0;
    assign memhint[6509] = 1'd0;
    assign memhint[6510] = 1'd0;
    assign memhint[6511] = 1'd0;
    assign memhint[6512] = 1'd0;
    assign memhint[6513] = 1'd0;
    assign memhint[6514] = 1'd0;
    assign memhint[6515] = 1'd0;
    assign memhint[6516] = 1'd0;
    assign memhint[6517] = 1'd0;
    assign memhint[6518] = 1'd0;
    assign memhint[6519] = 1'd0;
    assign memhint[6520] = 1'd0;
    assign memhint[6521] = 1'd0;
    assign memhint[6522] = 1'd0;
    assign memhint[6523] = 1'd1;
    assign memhint[6524] = 1'd1;
    assign memhint[6525] = 1'd0;
    assign memhint[6526] = 1'd0;
    assign memhint[6527] = 1'd0;
    assign memhint[6528] = 1'd0;
    assign memhint[6529] = 1'd0;
    assign memhint[6530] = 1'd0;
    assign memhint[6531] = 1'd0;
    assign memhint[6532] = 1'd1;
    assign memhint[6533] = 1'd1;
    assign memhint[6534] = 1'd0;
    assign memhint[6535] = 1'd0;
    assign memhint[6536] = 1'd0;
    assign memhint[6537] = 1'd0;
    assign memhint[6538] = 1'd0;
    assign memhint[6539] = 1'd0;
    assign memhint[6540] = 1'd0;
    assign memhint[6541] = 1'd0;
    assign memhint[6542] = 1'd0;
    assign memhint[6543] = 1'd0;
    assign memhint[6544] = 1'd0;
    assign memhint[6545] = 1'd1;
    assign memhint[6546] = 1'd1;
    assign memhint[6547] = 1'd0;
    assign memhint[6548] = 1'd1;
    assign memhint[6549] = 1'd1;
    assign memhint[6550] = 1'd0;
    assign memhint[6551] = 1'd0;
    assign memhint[6552] = 1'd0;
    assign memhint[6553] = 1'd0;
    assign memhint[6554] = 1'd0;
    assign memhint[6555] = 1'd0;
    assign memhint[6556] = 1'd0;
    assign memhint[6557] = 1'd1;
    assign memhint[6558] = 1'd1;
    assign memhint[6559] = 1'd0;
    assign memhint[6560] = 1'd0;
    assign memhint[6561] = 1'd0;
    assign memhint[6562] = 1'd0;
    assign memhint[6563] = 1'd0;
    assign memhint[6564] = 1'd0;
    assign memhint[6565] = 1'd0;
    assign memhint[6566] = 1'd0;
    assign memhint[6567] = 1'd0;
    assign memhint[6568] = 1'd0;
    assign memhint[6569] = 1'd0;
    assign memhint[6570] = 1'd0;
    assign memhint[6571] = 1'd0;
    assign memhint[6572] = 1'd0;
    assign memhint[6573] = 1'd0;
    assign memhint[6574] = 1'd0;
    assign memhint[6575] = 1'd0;
    assign memhint[6576] = 1'd1;
    assign memhint[6577] = 1'd1;
    assign memhint[6578] = 1'd0;
    assign memhint[6579] = 1'd0;
    assign memhint[6580] = 1'd0;
    assign memhint[6581] = 1'd0;
    assign memhint[6582] = 1'd0;
    assign memhint[6583] = 1'd0;
    assign memhint[6584] = 1'd0;
    assign memhint[6585] = 1'd0;
    assign memhint[6586] = 1'd0;
    assign memhint[6587] = 1'd0;
    assign memhint[6588] = 1'd0;
    assign memhint[6589] = 1'd0;
    assign memhint[6590] = 1'd0;
    assign memhint[6591] = 1'd0;
    assign memhint[6592] = 1'd0;
    assign memhint[6593] = 1'd0;
    assign memhint[6594] = 1'd0;
    assign memhint[6595] = 1'd1;
    assign memhint[6596] = 1'd1;
    assign memhint[6597] = 1'd0;
    assign memhint[6598] = 1'd0;
    assign memhint[6599] = 1'd0;
    assign memhint[6600] = 1'd0;
    assign memhint[6601] = 1'd0;
    assign memhint[6602] = 1'd0;
    assign memhint[6603] = 1'd0;
    assign memhint[6604] = 1'd0;
    assign memhint[6605] = 1'd0;
    assign memhint[6606] = 1'd0;
    assign memhint[6607] = 1'd1;
    assign memhint[6608] = 1'd1;
    assign memhint[6609] = 1'd0;
    assign memhint[6610] = 1'd0;
    assign memhint[6611] = 1'd0;
    assign memhint[6612] = 1'd0;
    assign memhint[6613] = 1'd0;
    assign memhint[6614] = 1'd0;
    assign memhint[6615] = 1'd0;
    assign memhint[6616] = 1'd0;
    assign memhint[6617] = 1'd0;
    assign memhint[6618] = 1'd0;
    assign memhint[6619] = 1'd0;
    assign memhint[6620] = 1'd0;
    assign memhint[6621] = 1'd0;
    assign memhint[6622] = 1'd0;
    assign memhint[6623] = 1'd0;
    assign memhint[6624] = 1'd0;
    assign memhint[6625] = 1'd1;
    assign memhint[6626] = 1'd1;
    assign memhint[6627] = 1'd0;
    assign memhint[6628] = 1'd0;
    assign memhint[6629] = 1'd0;
    assign memhint[6630] = 1'd0;
    assign memhint[6631] = 1'd0;
    assign memhint[6632] = 1'd0;
    assign memhint[6633] = 1'd0;
    assign memhint[6634] = 1'd0;
    assign memhint[6635] = 1'd0;
    assign memhint[6636] = 1'd0;
    assign memhint[6637] = 1'd0;
    assign memhint[6638] = 1'd0;
    assign memhint[6639] = 1'd0;
    assign memhint[6640] = 1'd0;
    assign memhint[6641] = 1'd0;
    assign memhint[6642] = 1'd0;
    assign memhint[6643] = 1'd1;
    assign memhint[6644] = 1'd1;
    assign memhint[6645] = 1'd0;
    assign memhint[6646] = 1'd0;
    assign memhint[6647] = 1'd0;
    assign memhint[6648] = 1'd0;
    assign memhint[6649] = 1'd0;
    assign memhint[6650] = 1'd0;
    assign memhint[6651] = 1'd0;
    assign memhint[6652] = 1'd0;
    assign memhint[6653] = 1'd0;
    assign memhint[6654] = 1'd0;
    assign memhint[6655] = 1'd0;
    assign memhint[6656] = 1'd0;
    assign memhint[6657] = 1'd0;
    assign memhint[6658] = 1'd0;
    assign memhint[6659] = 1'd0;
    assign memhint[6660] = 1'd0;
    assign memhint[6661] = 1'd0;
    assign memhint[6662] = 1'd1;
    assign memhint[6663] = 1'd1;
    assign memhint[6664] = 1'd0;
    assign memhint[6665] = 1'd0;
    assign memhint[6666] = 1'd0;
    assign memhint[6667] = 1'd0;
    assign memhint[6668] = 1'd0;
    assign memhint[6669] = 1'd0;
    assign memhint[6670] = 1'd0;
    assign memhint[6671] = 1'd0;
    assign memhint[6672] = 1'd0;
    assign memhint[6673] = 1'd0;
    assign memhint[6674] = 1'd0;
    assign memhint[6675] = 1'd0;
    assign memhint[6676] = 1'd0;
    assign memhint[6677] = 1'd1;
    assign memhint[6678] = 1'd1;
    assign memhint[6679] = 1'd1;
    assign memhint[6680] = 1'd0;
    assign memhint[6681] = 1'd0;
    assign memhint[6682] = 1'd0;
    assign memhint[6683] = 1'd0;
    assign memhint[6684] = 1'd0;
    assign memhint[6685] = 1'd0;
    assign memhint[6686] = 1'd0;
    assign memhint[6687] = 1'd0;
    assign memhint[6688] = 1'd0;
    assign memhint[6689] = 1'd0;
    assign memhint[6690] = 1'd0;
    assign memhint[6691] = 1'd0;
    assign memhint[6692] = 1'd1;
    assign memhint[6693] = 1'd1;
    assign memhint[6694] = 1'd0;
    assign memhint[6695] = 1'd0;
    assign memhint[6696] = 1'd0;
    assign memhint[6697] = 1'd0;
    assign memhint[6698] = 1'd0;
    assign memhint[6699] = 1'd0;
    assign memhint[6700] = 1'd0;
    assign memhint[6701] = 1'd0;
    assign memhint[6702] = 1'd0;
    assign memhint[6703] = 1'd0;
    assign memhint[6704] = 1'd0;
    assign memhint[6705] = 1'd1;
    assign memhint[6706] = 1'd1;
    assign memhint[6707] = 1'd0;
    assign memhint[6708] = 1'd0;
    assign memhint[6709] = 1'd0;
    assign memhint[6710] = 1'd0;
    assign memhint[6711] = 1'd0;
    assign memhint[6712] = 1'd0;
    assign memhint[6713] = 1'd0;
    assign memhint[6714] = 1'd1;
    assign memhint[6715] = 1'd1;
    assign memhint[6716] = 1'd1;
    assign memhint[6717] = 1'd0;
    assign memhint[6718] = 1'd0;
    assign memhint[6719] = 1'd0;
    assign memhint[6720] = 1'd0;
    assign memhint[6721] = 1'd0;
    assign memhint[6722] = 1'd0;
    assign memhint[6723] = 1'd0;
    assign memhint[6724] = 1'd0;
    assign memhint[6725] = 1'd1;
    assign memhint[6726] = 1'd1;
    assign memhint[6727] = 1'd0;
    assign memhint[6728] = 1'd0;
    assign memhint[6729] = 1'd0;
    assign memhint[6730] = 1'd0;
    assign memhint[6731] = 1'd0;
    assign memhint[6732] = 1'd1;
    assign memhint[6733] = 1'd1;
    assign memhint[6734] = 1'd0;
    assign memhint[6735] = 1'd0;
    assign memhint[6736] = 1'd0;
    assign memhint[6737] = 1'd0;
    assign memhint[6738] = 1'd0;
    assign memhint[6739] = 1'd0;
    assign memhint[6740] = 1'd0;
    assign memhint[6741] = 1'd0;
    assign memhint[6742] = 1'd0;
    assign memhint[6743] = 1'd0;
    assign memhint[6744] = 1'd0;
    assign memhint[6745] = 1'd0;
    assign memhint[6746] = 1'd0;
    assign memhint[6747] = 1'd0;
    assign memhint[6748] = 1'd0;
    assign memhint[6749] = 1'd1;
    assign memhint[6750] = 1'd1;
    assign memhint[6751] = 1'd0;
    assign memhint[6752] = 1'd0;
    assign memhint[6753] = 1'd0;
    assign memhint[6754] = 1'd0;
    assign memhint[6755] = 1'd0;
    assign memhint[6756] = 1'd0;
    assign memhint[6757] = 1'd0;
    assign memhint[6758] = 1'd0;
    assign memhint[6759] = 1'd0;
    assign memhint[6760] = 1'd0;
    assign memhint[6761] = 1'd0;
    assign memhint[6762] = 1'd0;
    assign memhint[6763] = 1'd0;
    assign memhint[6764] = 1'd1;
    assign memhint[6765] = 1'd1;
    assign memhint[6766] = 1'd0;
    assign memhint[6767] = 1'd0;
    assign memhint[6768] = 1'd0;
    assign memhint[6769] = 1'd0;
    assign memhint[6770] = 1'd0;
    assign memhint[6771] = 1'd0;
    assign memhint[6772] = 1'd0;
    assign memhint[6773] = 1'd0;
    assign memhint[6774] = 1'd0;
    assign memhint[6775] = 1'd0;
    assign memhint[6776] = 1'd0;
    assign memhint[6777] = 1'd0;
    assign memhint[6778] = 1'd0;
    assign memhint[6779] = 1'd0;
    assign memhint[6780] = 1'd0;
    assign memhint[6781] = 1'd0;
    assign memhint[6782] = 1'd1;
    assign memhint[6783] = 1'd1;
    assign memhint[6784] = 1'd1;
    assign memhint[6785] = 1'd0;
    assign memhint[6786] = 1'd0;
    assign memhint[6787] = 1'd0;
    assign memhint[6788] = 1'd0;
    assign memhint[6789] = 1'd0;
    assign memhint[6790] = 1'd0;
    assign memhint[6791] = 1'd0;
    assign memhint[6792] = 1'd0;
    assign memhint[6793] = 1'd0;
    assign memhint[6794] = 1'd0;
    assign memhint[6795] = 1'd0;
    assign memhint[6796] = 1'd0;
    assign memhint[6797] = 1'd0;
    assign memhint[6798] = 1'd0;
    assign memhint[6799] = 1'd1;
    assign memhint[6800] = 1'd1;
    assign memhint[6801] = 1'd1;
    assign memhint[6802] = 1'd0;
    assign memhint[6803] = 1'd0;
    assign memhint[6804] = 1'd0;
    assign memhint[6805] = 1'd0;
    assign memhint[6806] = 1'd0;
    assign memhint[6807] = 1'd0;
    assign memhint[6808] = 1'd0;
    assign memhint[6809] = 1'd1;
    assign memhint[6810] = 1'd1;
    assign memhint[6811] = 1'd0;
    assign memhint[6812] = 1'd0;
    assign memhint[6813] = 1'd0;
    assign memhint[6814] = 1'd0;
    assign memhint[6815] = 1'd0;
    assign memhint[6816] = 1'd0;
    assign memhint[6817] = 1'd0;
    assign memhint[6818] = 1'd0;
    assign memhint[6819] = 1'd0;
    assign memhint[6820] = 1'd0;
    assign memhint[6821] = 1'd0;
    assign memhint[6822] = 1'd0;
    assign memhint[6823] = 1'd0;
    assign memhint[6824] = 1'd0;
    assign memhint[6825] = 1'd0;
    assign memhint[6826] = 1'd0;
    assign memhint[6827] = 1'd0;
    assign memhint[6828] = 1'd0;
    assign memhint[6829] = 1'd1;
    assign memhint[6830] = 1'd1;
    assign memhint[6831] = 1'd0;
    assign memhint[6832] = 1'd0;
    assign memhint[6833] = 1'd0;
    assign memhint[6834] = 1'd0;
    assign memhint[6835] = 1'd0;
    assign memhint[6836] = 1'd0;
    assign memhint[6837] = 1'd0;
    assign memhint[6838] = 1'd0;
    assign memhint[6839] = 1'd0;
    assign memhint[6840] = 1'd0;
    assign memhint[6841] = 1'd0;
    assign memhint[6842] = 1'd0;
    assign memhint[6843] = 1'd0;
    assign memhint[6844] = 1'd1;
    assign memhint[6845] = 1'd1;
    assign memhint[6846] = 1'd0;
    assign memhint[6847] = 1'd0;
    assign memhint[6848] = 1'd0;
    assign memhint[6849] = 1'd0;
    assign memhint[6850] = 1'd0;
    assign memhint[6851] = 1'd0;
    assign memhint[6852] = 1'd0;
    assign memhint[6853] = 1'd0;
    assign memhint[6854] = 1'd0;
    assign memhint[6855] = 1'd0;
    assign memhint[6856] = 1'd0;
    assign memhint[6857] = 1'd0;
    assign memhint[6858] = 1'd0;
    assign memhint[6859] = 1'd1;
    assign memhint[6860] = 1'd1;
    assign memhint[6861] = 1'd1;
    assign memhint[6862] = 1'd0;
    assign memhint[6863] = 1'd0;
    assign memhint[6864] = 1'd0;
    assign memhint[6865] = 1'd0;
    assign memhint[6866] = 1'd0;
    assign memhint[6867] = 1'd0;
    assign memhint[6868] = 1'd0;
    assign memhint[6869] = 1'd0;
    assign memhint[6870] = 1'd1;
    assign memhint[6871] = 1'd1;
    assign memhint[6872] = 1'd0;
    assign memhint[6873] = 1'd0;
    assign memhint[6874] = 1'd0;
    assign memhint[6875] = 1'd0;
    assign memhint[6876] = 1'd0;
    assign memhint[6877] = 1'd0;
    assign memhint[6878] = 1'd1;
    assign memhint[6879] = 1'd1;
    assign memhint[6880] = 1'd1;
    assign memhint[6881] = 1'd0;
    assign memhint[6882] = 1'd0;
    assign memhint[6883] = 1'd0;
    assign memhint[6884] = 1'd0;
    assign memhint[6885] = 1'd0;
    assign memhint[6886] = 1'd0;
    assign memhint[6887] = 1'd0;
    assign memhint[6888] = 1'd0;
    assign memhint[6889] = 1'd0;
    assign memhint[6890] = 1'd0;
    assign memhint[6891] = 1'd0;
    assign memhint[6892] = 1'd0;
    assign memhint[6893] = 1'd0;
    assign memhint[6894] = 1'd0;
    assign memhint[6895] = 1'd1;
    assign memhint[6896] = 1'd1;
    assign memhint[6897] = 1'd1;
    assign memhint[6898] = 1'd0;
    assign memhint[6899] = 1'd0;
    assign memhint[6900] = 1'd0;
    assign memhint[6901] = 1'd0;
    assign memhint[6902] = 1'd0;
    assign memhint[6903] = 1'd0;
    assign memhint[6904] = 1'd0;
    assign memhint[6905] = 1'd1;
    assign memhint[6906] = 1'd1;
    assign memhint[6907] = 1'd0;
    assign memhint[6908] = 1'd0;
    assign memhint[6909] = 1'd0;
    assign memhint[6910] = 1'd0;
    assign memhint[6911] = 1'd0;
    assign memhint[6912] = 1'd0;
    assign memhint[6913] = 1'd0;
    assign memhint[6914] = 1'd0;
    assign memhint[6915] = 1'd0;
    assign memhint[6916] = 1'd0;
    assign memhint[6917] = 1'd0;
    assign memhint[6918] = 1'd0;
    assign memhint[6919] = 1'd1;
    assign memhint[6920] = 1'd1;
    assign memhint[6921] = 1'd1;
    assign memhint[6922] = 1'd1;
    assign memhint[6923] = 1'd0;
    assign memhint[6924] = 1'd0;
    assign memhint[6925] = 1'd0;
    assign memhint[6926] = 1'd0;
    assign memhint[6927] = 1'd0;
    assign memhint[6928] = 1'd0;
    assign memhint[6929] = 1'd0;
    assign memhint[6930] = 1'd1;
    assign memhint[6931] = 1'd1;
    assign memhint[6932] = 1'd1;
    assign memhint[6933] = 1'd0;
    assign memhint[6934] = 1'd0;
    assign memhint[6935] = 1'd0;
    assign memhint[6936] = 1'd0;
    assign memhint[6937] = 1'd0;
    assign memhint[6938] = 1'd0;
    assign memhint[6939] = 1'd0;
    assign memhint[6940] = 1'd0;
    assign memhint[6941] = 1'd0;
    assign memhint[6942] = 1'd0;
    assign memhint[6943] = 1'd0;
    assign memhint[6944] = 1'd0;
    assign memhint[6945] = 1'd0;
    assign memhint[6946] = 1'd0;
    assign memhint[6947] = 1'd0;
    assign memhint[6948] = 1'd1;
    assign memhint[6949] = 1'd1;
    assign memhint[6950] = 1'd0;
    assign memhint[6951] = 1'd0;
    assign memhint[6952] = 1'd0;
    assign memhint[6953] = 1'd0;
    assign memhint[6954] = 1'd0;
    assign memhint[6955] = 1'd0;
    assign memhint[6956] = 1'd0;
    assign memhint[6957] = 1'd0;
    assign memhint[6958] = 1'd0;
    assign memhint[6959] = 1'd0;
    assign memhint[6960] = 1'd0;
    assign memhint[6961] = 1'd0;
    assign memhint[6962] = 1'd0;
    assign memhint[6963] = 1'd0;
    assign memhint[6964] = 1'd0;
    assign memhint[6965] = 1'd0;
    assign memhint[6966] = 1'd0;
    assign memhint[6967] = 1'd0;
    assign memhint[6968] = 1'd1;
    assign memhint[6969] = 1'd1;
    assign memhint[6970] = 1'd0;
    assign memhint[6971] = 1'd0;
    assign memhint[6972] = 1'd0;
    assign memhint[6973] = 1'd0;
    assign memhint[6974] = 1'd0;
    assign memhint[6975] = 1'd0;
    assign memhint[6976] = 1'd0;
    assign memhint[6977] = 1'd0;
    assign memhint[6978] = 1'd0;
    assign memhint[6979] = 1'd0;
    assign memhint[6980] = 1'd1;
    assign memhint[6981] = 1'd1;
    assign memhint[6982] = 1'd1;
    assign memhint[6983] = 1'd0;
    assign memhint[6984] = 1'd0;
    assign memhint[6985] = 1'd0;
    assign memhint[6986] = 1'd0;
    assign memhint[6987] = 1'd0;
    assign memhint[6988] = 1'd0;
    assign memhint[6989] = 1'd0;
    assign memhint[6990] = 1'd0;
    assign memhint[6991] = 1'd0;
    assign memhint[6992] = 1'd0;
    assign memhint[6993] = 1'd0;
    assign memhint[6994] = 1'd0;
    assign memhint[6995] = 1'd0;
    assign memhint[6996] = 1'd0;
    assign memhint[6997] = 1'd1;
    assign memhint[6998] = 1'd1;
    assign memhint[6999] = 1'd1;
    assign memhint[7000] = 1'd0;
    assign memhint[7001] = 1'd0;
    assign memhint[7002] = 1'd0;
    assign memhint[7003] = 1'd0;
    assign memhint[7004] = 1'd0;
    assign memhint[7005] = 1'd0;
    assign memhint[7006] = 1'd0;
    assign memhint[7007] = 1'd0;
    assign memhint[7008] = 1'd0;
    assign memhint[7009] = 1'd0;
    assign memhint[7010] = 1'd0;
    assign memhint[7011] = 1'd0;
    assign memhint[7012] = 1'd0;
    assign memhint[7013] = 1'd0;
    assign memhint[7014] = 1'd0;
    assign memhint[7015] = 1'd0;
    assign memhint[7016] = 1'd1;
    assign memhint[7017] = 1'd1;
    assign memhint[7018] = 1'd0;
    assign memhint[7019] = 1'd0;
    assign memhint[7020] = 1'd0;
    assign memhint[7021] = 1'd0;
    assign memhint[7022] = 1'd0;
    assign memhint[7023] = 1'd0;
    assign memhint[7024] = 1'd0;
    assign memhint[7025] = 1'd0;
    assign memhint[7026] = 1'd0;
    assign memhint[7027] = 1'd0;
    assign memhint[7028] = 1'd0;
    assign memhint[7029] = 1'd0;
    assign memhint[7030] = 1'd0;
    assign memhint[7031] = 1'd0;
    assign memhint[7032] = 1'd0;
    assign memhint[7033] = 1'd0;
    assign memhint[7034] = 1'd0;
    assign memhint[7035] = 1'd1;
    assign memhint[7036] = 1'd1;
    assign memhint[7037] = 1'd0;
    assign memhint[7038] = 1'd0;
    assign memhint[7039] = 1'd0;
    assign memhint[7040] = 1'd0;
    assign memhint[7041] = 1'd0;
    assign memhint[7042] = 1'd0;
    assign memhint[7043] = 1'd0;
    assign memhint[7044] = 1'd0;
    assign memhint[7045] = 1'd0;
    assign memhint[7046] = 1'd0;
    assign memhint[7047] = 1'd0;
    assign memhint[7048] = 1'd0;
    assign memhint[7049] = 1'd0;
    assign memhint[7050] = 1'd1;
    assign memhint[7051] = 1'd1;
    assign memhint[7052] = 1'd0;
    assign memhint[7053] = 1'd0;
    assign memhint[7054] = 1'd0;
    assign memhint[7055] = 1'd0;
    assign memhint[7056] = 1'd0;
    assign memhint[7057] = 1'd0;
    assign memhint[7058] = 1'd0;
    assign memhint[7059] = 1'd0;
    assign memhint[7060] = 1'd0;
    assign memhint[7061] = 1'd0;
    assign memhint[7062] = 1'd0;
    assign memhint[7063] = 1'd0;
    assign memhint[7064] = 1'd0;
    assign memhint[7065] = 1'd1;
    assign memhint[7066] = 1'd1;
    assign memhint[7067] = 1'd0;
    assign memhint[7068] = 1'd0;
    assign memhint[7069] = 1'd0;
    assign memhint[7070] = 1'd0;
    assign memhint[7071] = 1'd0;
    assign memhint[7072] = 1'd0;
    assign memhint[7073] = 1'd0;
    assign memhint[7074] = 1'd0;
    assign memhint[7075] = 1'd0;
    assign memhint[7076] = 1'd0;
    assign memhint[7077] = 1'd0;
    assign memhint[7078] = 1'd1;
    assign memhint[7079] = 1'd1;
    assign memhint[7080] = 1'd0;
    assign memhint[7081] = 1'd0;
    assign memhint[7082] = 1'd0;
    assign memhint[7083] = 1'd0;
    assign memhint[7084] = 1'd0;
    assign memhint[7085] = 1'd0;
    assign memhint[7086] = 1'd0;
    assign memhint[7087] = 1'd0;
    assign memhint[7088] = 1'd1;
    assign memhint[7089] = 1'd1;
    assign memhint[7090] = 1'd1;
    assign memhint[7091] = 1'd0;
    assign memhint[7092] = 1'd0;
    assign memhint[7093] = 1'd0;
    assign memhint[7094] = 1'd0;
    assign memhint[7095] = 1'd0;
    assign memhint[7096] = 1'd0;
    assign memhint[7097] = 1'd1;
    assign memhint[7098] = 1'd1;
    assign memhint[7099] = 1'd0;
    assign memhint[7100] = 1'd0;
    assign memhint[7101] = 1'd0;
    assign memhint[7102] = 1'd0;
    assign memhint[7103] = 1'd0;
    assign memhint[7104] = 1'd0;
    assign memhint[7105] = 1'd1;
    assign memhint[7106] = 1'd1;
    assign memhint[7107] = 1'd0;
    assign memhint[7108] = 1'd0;
    assign memhint[7109] = 1'd0;
    assign memhint[7110] = 1'd0;
    assign memhint[7111] = 1'd0;
    assign memhint[7112] = 1'd0;
    assign memhint[7113] = 1'd0;
    assign memhint[7114] = 1'd0;
    assign memhint[7115] = 1'd0;
    assign memhint[7116] = 1'd0;
    assign memhint[7117] = 1'd0;
    assign memhint[7118] = 1'd0;
    assign memhint[7119] = 1'd0;
    assign memhint[7120] = 1'd0;
    assign memhint[7121] = 1'd0;
    assign memhint[7122] = 1'd1;
    assign memhint[7123] = 1'd1;
    assign memhint[7124] = 1'd0;
    assign memhint[7125] = 1'd0;
    assign memhint[7126] = 1'd0;
    assign memhint[7127] = 1'd0;
    assign memhint[7128] = 1'd0;
    assign memhint[7129] = 1'd0;
    assign memhint[7130] = 1'd0;
    assign memhint[7131] = 1'd0;
    assign memhint[7132] = 1'd0;
    assign memhint[7133] = 1'd0;
    assign memhint[7134] = 1'd0;
    assign memhint[7135] = 1'd0;
    assign memhint[7136] = 1'd0;
    assign memhint[7137] = 1'd1;
    assign memhint[7138] = 1'd1;
    assign memhint[7139] = 1'd0;
    assign memhint[7140] = 1'd0;
    assign memhint[7141] = 1'd0;
    assign memhint[7142] = 1'd0;
    assign memhint[7143] = 1'd0;
    assign memhint[7144] = 1'd0;
    assign memhint[7145] = 1'd0;
    assign memhint[7146] = 1'd0;
    assign memhint[7147] = 1'd0;
    assign memhint[7148] = 1'd0;
    assign memhint[7149] = 1'd0;
    assign memhint[7150] = 1'd0;
    assign memhint[7151] = 1'd0;
    assign memhint[7152] = 1'd0;
    assign memhint[7153] = 1'd0;
    assign memhint[7154] = 1'd0;
    assign memhint[7155] = 1'd0;
    assign memhint[7156] = 1'd1;
    assign memhint[7157] = 1'd1;
    assign memhint[7158] = 1'd1;
    assign memhint[7159] = 1'd0;
    assign memhint[7160] = 1'd0;
    assign memhint[7161] = 1'd0;
    assign memhint[7162] = 1'd0;
    assign memhint[7163] = 1'd0;
    assign memhint[7164] = 1'd0;
    assign memhint[7165] = 1'd0;
    assign memhint[7166] = 1'd0;
    assign memhint[7167] = 1'd0;
    assign memhint[7168] = 1'd0;
    assign memhint[7169] = 1'd0;
    assign memhint[7170] = 1'd1;
    assign memhint[7171] = 1'd1;
    assign memhint[7172] = 1'd1;
    assign memhint[7173] = 1'd1;
    assign memhint[7174] = 1'd0;
    assign memhint[7175] = 1'd0;
    assign memhint[7176] = 1'd0;
    assign memhint[7177] = 1'd0;
    assign memhint[7178] = 1'd0;
    assign memhint[7179] = 1'd0;
    assign memhint[7180] = 1'd0;
    assign memhint[7181] = 1'd0;
    assign memhint[7182] = 1'd1;
    assign memhint[7183] = 1'd1;
    assign memhint[7184] = 1'd0;
    assign memhint[7185] = 1'd0;
    assign memhint[7186] = 1'd0;
    assign memhint[7187] = 1'd0;
    assign memhint[7188] = 1'd0;
    assign memhint[7189] = 1'd0;
    assign memhint[7190] = 1'd0;
    assign memhint[7191] = 1'd0;
    assign memhint[7192] = 1'd0;
    assign memhint[7193] = 1'd0;
    assign memhint[7194] = 1'd0;
    assign memhint[7195] = 1'd0;
    assign memhint[7196] = 1'd0;
    assign memhint[7197] = 1'd0;
    assign memhint[7198] = 1'd0;
    assign memhint[7199] = 1'd0;
    assign memhint[7200] = 1'd0;
    assign memhint[7201] = 1'd0;
    assign memhint[7202] = 1'd1;
    assign memhint[7203] = 1'd1;
    assign memhint[7204] = 1'd0;
    assign memhint[7205] = 1'd0;
    assign memhint[7206] = 1'd0;
    assign memhint[7207] = 1'd0;
    assign memhint[7208] = 1'd0;
    assign memhint[7209] = 1'd0;
    assign memhint[7210] = 1'd0;
    assign memhint[7211] = 1'd0;
    assign memhint[7212] = 1'd0;
    assign memhint[7213] = 1'd0;
    assign memhint[7214] = 1'd0;
    assign memhint[7215] = 1'd0;
    assign memhint[7216] = 1'd0;
    assign memhint[7217] = 1'd1;
    assign memhint[7218] = 1'd1;
    assign memhint[7219] = 1'd0;
    assign memhint[7220] = 1'd0;
    assign memhint[7221] = 1'd0;
    assign memhint[7222] = 1'd0;
    assign memhint[7223] = 1'd0;
    assign memhint[7224] = 1'd0;
    assign memhint[7225] = 1'd0;
    assign memhint[7226] = 1'd0;
    assign memhint[7227] = 1'd0;
    assign memhint[7228] = 1'd0;
    assign memhint[7229] = 1'd0;
    assign memhint[7230] = 1'd0;
    assign memhint[7231] = 1'd0;
    assign memhint[7232] = 1'd0;
    assign memhint[7233] = 1'd1;
    assign memhint[7234] = 1'd1;
    assign memhint[7235] = 1'd1;
    assign memhint[7236] = 1'd0;
    assign memhint[7237] = 1'd0;
    assign memhint[7238] = 1'd0;
    assign memhint[7239] = 1'd0;
    assign memhint[7240] = 1'd0;
    assign memhint[7241] = 1'd0;
    assign memhint[7242] = 1'd1;
    assign memhint[7243] = 1'd1;
    assign memhint[7244] = 1'd0;
    assign memhint[7245] = 1'd0;
    assign memhint[7246] = 1'd0;
    assign memhint[7247] = 1'd0;
    assign memhint[7248] = 1'd0;
    assign memhint[7249] = 1'd0;
    assign memhint[7250] = 1'd0;
    assign memhint[7251] = 1'd0;
    assign memhint[7252] = 1'd1;
    assign memhint[7253] = 1'd1;
    assign memhint[7254] = 1'd1;
    assign memhint[7255] = 1'd1;
    assign memhint[7256] = 1'd0;
    assign memhint[7257] = 1'd0;
    assign memhint[7258] = 1'd0;
    assign memhint[7259] = 1'd0;
    assign memhint[7260] = 1'd0;
    assign memhint[7261] = 1'd0;
    assign memhint[7262] = 1'd0;
    assign memhint[7263] = 1'd0;
    assign memhint[7264] = 1'd0;
    assign memhint[7265] = 1'd0;
    assign memhint[7266] = 1'd1;
    assign memhint[7267] = 1'd1;
    assign memhint[7268] = 1'd1;
    assign memhint[7269] = 1'd1;
    assign memhint[7270] = 1'd0;
    assign memhint[7271] = 1'd0;
    assign memhint[7272] = 1'd0;
    assign memhint[7273] = 1'd0;
    assign memhint[7274] = 1'd0;
    assign memhint[7275] = 1'd0;
    assign memhint[7276] = 1'd0;
    assign memhint[7277] = 1'd0;
    assign memhint[7278] = 1'd1;
    assign memhint[7279] = 1'd1;
    assign memhint[7280] = 1'd0;
    assign memhint[7281] = 1'd0;
    assign memhint[7282] = 1'd0;
    assign memhint[7283] = 1'd0;
    assign memhint[7284] = 1'd0;
    assign memhint[7285] = 1'd0;
    assign memhint[7286] = 1'd0;
    assign memhint[7287] = 1'd0;
    assign memhint[7288] = 1'd0;
    assign memhint[7289] = 1'd0;
    assign memhint[7290] = 1'd0;
    assign memhint[7291] = 1'd0;
    assign memhint[7292] = 1'd0;
    assign memhint[7293] = 1'd1;
    assign memhint[7294] = 1'd1;
    assign memhint[7295] = 1'd1;
    assign memhint[7296] = 1'd0;
    assign memhint[7297] = 1'd0;
    assign memhint[7298] = 1'd0;
    assign memhint[7299] = 1'd0;
    assign memhint[7300] = 1'd0;
    assign memhint[7301] = 1'd0;
    assign memhint[7302] = 1'd0;
    assign memhint[7303] = 1'd0;
    assign memhint[7304] = 1'd1;
    assign memhint[7305] = 1'd1;
    assign memhint[7306] = 1'd1;
    assign memhint[7307] = 1'd1;
    assign memhint[7308] = 1'd0;
    assign memhint[7309] = 1'd0;
    assign memhint[7310] = 1'd0;
    assign memhint[7311] = 1'd0;
    assign memhint[7312] = 1'd0;
    assign memhint[7313] = 1'd0;
    assign memhint[7314] = 1'd0;
    assign memhint[7315] = 1'd0;
    assign memhint[7316] = 1'd0;
    assign memhint[7317] = 1'd0;
    assign memhint[7318] = 1'd0;
    assign memhint[7319] = 1'd1;
    assign memhint[7320] = 1'd1;
    assign memhint[7321] = 1'd1;
    assign memhint[7322] = 1'd0;
    assign memhint[7323] = 1'd0;
    assign memhint[7324] = 1'd0;
    assign memhint[7325] = 1'd0;
    assign memhint[7326] = 1'd0;
    assign memhint[7327] = 1'd0;
    assign memhint[7328] = 1'd0;
    assign memhint[7329] = 1'd0;
    assign memhint[7330] = 1'd0;
    assign memhint[7331] = 1'd0;
    assign memhint[7332] = 1'd0;
    assign memhint[7333] = 1'd0;
    assign memhint[7334] = 1'd0;
    assign memhint[7335] = 1'd0;
    assign memhint[7336] = 1'd0;
    assign memhint[7337] = 1'd0;
    assign memhint[7338] = 1'd0;
    assign memhint[7339] = 1'd0;
    assign memhint[7340] = 1'd0;
    assign memhint[7341] = 1'd1;
    assign memhint[7342] = 1'd1;
    assign memhint[7343] = 1'd0;
    assign memhint[7344] = 1'd0;
    assign memhint[7345] = 1'd0;
    assign memhint[7346] = 1'd0;
    assign memhint[7347] = 1'd0;
    assign memhint[7348] = 1'd0;
    assign memhint[7349] = 1'd0;
    assign memhint[7350] = 1'd0;
    assign memhint[7351] = 1'd0;
    assign memhint[7352] = 1'd0;
    assign memhint[7353] = 1'd0;
    assign memhint[7354] = 1'd1;
    assign memhint[7355] = 1'd1;
    assign memhint[7356] = 1'd1;
    assign memhint[7357] = 1'd1;
    assign memhint[7358] = 1'd0;
    assign memhint[7359] = 1'd0;
    assign memhint[7360] = 1'd0;
    assign memhint[7361] = 1'd0;
    assign memhint[7362] = 1'd0;
    assign memhint[7363] = 1'd0;
    assign memhint[7364] = 1'd0;
    assign memhint[7365] = 1'd0;
    assign memhint[7366] = 1'd0;
    assign memhint[7367] = 1'd0;
    assign memhint[7368] = 1'd1;
    assign memhint[7369] = 1'd1;
    assign memhint[7370] = 1'd1;
    assign memhint[7371] = 1'd1;
    assign memhint[7372] = 1'd0;
    assign memhint[7373] = 1'd0;
    assign memhint[7374] = 1'd0;
    assign memhint[7375] = 1'd0;
    assign memhint[7376] = 1'd0;
    assign memhint[7377] = 1'd0;
    assign memhint[7378] = 1'd0;
    assign memhint[7379] = 1'd0;
    assign memhint[7380] = 1'd0;
    assign memhint[7381] = 1'd0;
    assign memhint[7382] = 1'd0;
    assign memhint[7383] = 1'd0;
    assign memhint[7384] = 1'd0;
    assign memhint[7385] = 1'd0;
    assign memhint[7386] = 1'd0;
    assign memhint[7387] = 1'd0;
    assign memhint[7388] = 1'd0;
    assign memhint[7389] = 1'd1;
    assign memhint[7390] = 1'd1;
    assign memhint[7391] = 1'd0;
    assign memhint[7392] = 1'd0;
    assign memhint[7393] = 1'd0;
    assign memhint[7394] = 1'd0;
    assign memhint[7395] = 1'd0;
    assign memhint[7396] = 1'd0;
    assign memhint[7397] = 1'd0;
    assign memhint[7398] = 1'd0;
    assign memhint[7399] = 1'd0;
    assign memhint[7400] = 1'd0;
    assign memhint[7401] = 1'd0;
    assign memhint[7402] = 1'd0;
    assign memhint[7403] = 1'd0;
    assign memhint[7404] = 1'd0;
    assign memhint[7405] = 1'd0;
    assign memhint[7406] = 1'd0;
    assign memhint[7407] = 1'd0;
    assign memhint[7408] = 1'd1;
    assign memhint[7409] = 1'd1;
    assign memhint[7410] = 1'd0;
    assign memhint[7411] = 1'd0;
    assign memhint[7412] = 1'd0;
    assign memhint[7413] = 1'd0;
    assign memhint[7414] = 1'd0;
    assign memhint[7415] = 1'd0;
    assign memhint[7416] = 1'd0;
    assign memhint[7417] = 1'd0;
    assign memhint[7418] = 1'd0;
    assign memhint[7419] = 1'd0;
    assign memhint[7420] = 1'd0;
    assign memhint[7421] = 1'd0;
    assign memhint[7422] = 1'd0;
    assign memhint[7423] = 1'd1;
    assign memhint[7424] = 1'd1;
    assign memhint[7425] = 1'd0;
    assign memhint[7426] = 1'd0;
    assign memhint[7427] = 1'd0;
    assign memhint[7428] = 1'd0;
    assign memhint[7429] = 1'd0;
    assign memhint[7430] = 1'd0;
    assign memhint[7431] = 1'd0;
    assign memhint[7432] = 1'd0;
    assign memhint[7433] = 1'd0;
    assign memhint[7434] = 1'd0;
    assign memhint[7435] = 1'd0;
    assign memhint[7436] = 1'd0;
    assign memhint[7437] = 1'd0;
    assign memhint[7438] = 1'd1;
    assign memhint[7439] = 1'd1;
    assign memhint[7440] = 1'd0;
    assign memhint[7441] = 1'd0;
    assign memhint[7442] = 1'd0;
    assign memhint[7443] = 1'd0;
    assign memhint[7444] = 1'd0;
    assign memhint[7445] = 1'd0;
    assign memhint[7446] = 1'd0;
    assign memhint[7447] = 1'd0;
    assign memhint[7448] = 1'd0;
    assign memhint[7449] = 1'd0;
    assign memhint[7450] = 1'd0;
    assign memhint[7451] = 1'd1;
    assign memhint[7452] = 1'd1;
    assign memhint[7453] = 1'd0;
    assign memhint[7454] = 1'd0;
    assign memhint[7455] = 1'd0;
    assign memhint[7456] = 1'd0;
    assign memhint[7457] = 1'd0;
    assign memhint[7458] = 1'd0;
    assign memhint[7459] = 1'd0;
    assign memhint[7460] = 1'd0;
    assign memhint[7461] = 1'd0;
    assign memhint[7462] = 1'd1;
    assign memhint[7463] = 1'd1;
    assign memhint[7464] = 1'd1;
    assign memhint[7465] = 1'd0;
    assign memhint[7466] = 1'd0;
    assign memhint[7467] = 1'd0;
    assign memhint[7468] = 1'd0;
    assign memhint[7469] = 1'd1;
    assign memhint[7470] = 1'd1;
    assign memhint[7471] = 1'd1;
    assign memhint[7472] = 1'd0;
    assign memhint[7473] = 1'd0;
    assign memhint[7474] = 1'd0;
    assign memhint[7475] = 1'd0;
    assign memhint[7476] = 1'd0;
    assign memhint[7477] = 1'd0;
    assign memhint[7478] = 1'd1;
    assign memhint[7479] = 1'd1;
    assign memhint[7480] = 1'd0;
    assign memhint[7481] = 1'd0;
    assign memhint[7482] = 1'd0;
    assign memhint[7483] = 1'd0;
    assign memhint[7484] = 1'd0;
    assign memhint[7485] = 1'd0;
    assign memhint[7486] = 1'd0;
    assign memhint[7487] = 1'd0;
    assign memhint[7488] = 1'd0;
    assign memhint[7489] = 1'd0;
    assign memhint[7490] = 1'd0;
    assign memhint[7491] = 1'd0;
    assign memhint[7492] = 1'd0;
    assign memhint[7493] = 1'd0;
    assign memhint[7494] = 1'd0;
    assign memhint[7495] = 1'd1;
    assign memhint[7496] = 1'd1;
    assign memhint[7497] = 1'd0;
    assign memhint[7498] = 1'd0;
    assign memhint[7499] = 1'd0;
    assign memhint[7500] = 1'd0;
    assign memhint[7501] = 1'd0;
    assign memhint[7502] = 1'd0;
    assign memhint[7503] = 1'd0;
    assign memhint[7504] = 1'd0;
    assign memhint[7505] = 1'd0;
    assign memhint[7506] = 1'd0;
    assign memhint[7507] = 1'd0;
    assign memhint[7508] = 1'd0;
    assign memhint[7509] = 1'd0;
    assign memhint[7510] = 1'd1;
    assign memhint[7511] = 1'd1;
    assign memhint[7512] = 1'd0;
    assign memhint[7513] = 1'd0;
    assign memhint[7514] = 1'd0;
    assign memhint[7515] = 1'd0;
    assign memhint[7516] = 1'd0;
    assign memhint[7517] = 1'd0;
    assign memhint[7518] = 1'd0;
    assign memhint[7519] = 1'd0;
    assign memhint[7520] = 1'd0;
    assign memhint[7521] = 1'd0;
    assign memhint[7522] = 1'd0;
    assign memhint[7523] = 1'd0;
    assign memhint[7524] = 1'd0;
    assign memhint[7525] = 1'd0;
    assign memhint[7526] = 1'd0;
    assign memhint[7527] = 1'd0;
    assign memhint[7528] = 1'd0;
    assign memhint[7529] = 1'd0;
    assign memhint[7530] = 1'd1;
    assign memhint[7531] = 1'd1;
    assign memhint[7532] = 1'd1;
    assign memhint[7533] = 1'd1;
    assign memhint[7534] = 1'd1;
    assign memhint[7535] = 1'd0;
    assign memhint[7536] = 1'd0;
    assign memhint[7537] = 1'd0;
    assign memhint[7538] = 1'd0;
    assign memhint[7539] = 1'd0;
    assign memhint[7540] = 1'd0;
    assign memhint[7541] = 1'd1;
    assign memhint[7542] = 1'd1;
    assign memhint[7543] = 1'd1;
    assign memhint[7544] = 1'd1;
    assign memhint[7545] = 1'd1;
    assign memhint[7546] = 1'd0;
    assign memhint[7547] = 1'd0;
    assign memhint[7548] = 1'd0;
    assign memhint[7549] = 1'd0;
    assign memhint[7550] = 1'd0;
    assign memhint[7551] = 1'd0;
    assign memhint[7552] = 1'd0;
    assign memhint[7553] = 1'd0;
    assign memhint[7554] = 1'd0;
    assign memhint[7555] = 1'd1;
    assign memhint[7556] = 1'd1;
    assign memhint[7557] = 1'd0;
    assign memhint[7558] = 1'd0;
    assign memhint[7559] = 1'd0;
    assign memhint[7560] = 1'd0;
    assign memhint[7561] = 1'd0;
    assign memhint[7562] = 1'd0;
    assign memhint[7563] = 1'd0;
    assign memhint[7564] = 1'd0;
    assign memhint[7565] = 1'd0;
    assign memhint[7566] = 1'd0;
    assign memhint[7567] = 1'd0;
    assign memhint[7568] = 1'd0;
    assign memhint[7569] = 1'd0;
    assign memhint[7570] = 1'd0;
    assign memhint[7571] = 1'd0;
    assign memhint[7572] = 1'd0;
    assign memhint[7573] = 1'd0;
    assign memhint[7574] = 1'd1;
    assign memhint[7575] = 1'd1;
    assign memhint[7576] = 1'd0;
    assign memhint[7577] = 1'd0;
    assign memhint[7578] = 1'd0;
    assign memhint[7579] = 1'd0;
    assign memhint[7580] = 1'd0;
    assign memhint[7581] = 1'd0;
    assign memhint[7582] = 1'd0;
    assign memhint[7583] = 1'd0;
    assign memhint[7584] = 1'd0;
    assign memhint[7585] = 1'd0;
    assign memhint[7586] = 1'd0;
    assign memhint[7587] = 1'd0;
    assign memhint[7588] = 1'd0;
    assign memhint[7589] = 1'd0;
    assign memhint[7590] = 1'd0;
    assign memhint[7591] = 1'd1;
    assign memhint[7592] = 1'd1;
    assign memhint[7593] = 1'd0;
    assign memhint[7594] = 1'd0;
    assign memhint[7595] = 1'd0;
    assign memhint[7596] = 1'd0;
    assign memhint[7597] = 1'd0;
    assign memhint[7598] = 1'd0;
    assign memhint[7599] = 1'd0;
    assign memhint[7600] = 1'd0;
    assign memhint[7601] = 1'd0;
    assign memhint[7602] = 1'd0;
    assign memhint[7603] = 1'd0;
    assign memhint[7604] = 1'd0;
    assign memhint[7605] = 1'd0;
    assign memhint[7606] = 1'd0;
    assign memhint[7607] = 1'd1;
    assign memhint[7608] = 1'd1;
    assign memhint[7609] = 1'd1;
    assign memhint[7610] = 1'd0;
    assign memhint[7611] = 1'd0;
    assign memhint[7612] = 1'd0;
    assign memhint[7613] = 1'd0;
    assign memhint[7614] = 1'd1;
    assign memhint[7615] = 1'd1;
    assign memhint[7616] = 1'd1;
    assign memhint[7617] = 1'd0;
    assign memhint[7618] = 1'd0;
    assign memhint[7619] = 1'd0;
    assign memhint[7620] = 1'd0;
    assign memhint[7621] = 1'd0;
    assign memhint[7622] = 1'd0;
    assign memhint[7623] = 1'd0;
    assign memhint[7624] = 1'd0;
    assign memhint[7625] = 1'd0;
    assign memhint[7626] = 1'd1;
    assign memhint[7627] = 1'd1;
    assign memhint[7628] = 1'd1;
    assign memhint[7629] = 1'd1;
    assign memhint[7630] = 1'd1;
    assign memhint[7631] = 1'd0;
    assign memhint[7632] = 1'd0;
    assign memhint[7633] = 1'd0;
    assign memhint[7634] = 1'd0;
    assign memhint[7635] = 1'd0;
    assign memhint[7636] = 1'd0;
    assign memhint[7637] = 1'd1;
    assign memhint[7638] = 1'd1;
    assign memhint[7639] = 1'd1;
    assign memhint[7640] = 1'd1;
    assign memhint[7641] = 1'd1;
    assign memhint[7642] = 1'd0;
    assign memhint[7643] = 1'd0;
    assign memhint[7644] = 1'd0;
    assign memhint[7645] = 1'd0;
    assign memhint[7646] = 1'd0;
    assign memhint[7647] = 1'd0;
    assign memhint[7648] = 1'd0;
    assign memhint[7649] = 1'd0;
    assign memhint[7650] = 1'd0;
    assign memhint[7651] = 1'd1;
    assign memhint[7652] = 1'd1;
    assign memhint[7653] = 1'd0;
    assign memhint[7654] = 1'd0;
    assign memhint[7655] = 1'd0;
    assign memhint[7656] = 1'd0;
    assign memhint[7657] = 1'd0;
    assign memhint[7658] = 1'd0;
    assign memhint[7659] = 1'd0;
    assign memhint[7660] = 1'd0;
    assign memhint[7661] = 1'd0;
    assign memhint[7662] = 1'd0;
    assign memhint[7663] = 1'd0;
    assign memhint[7664] = 1'd0;
    assign memhint[7665] = 1'd0;
    assign memhint[7666] = 1'd1;
    assign memhint[7667] = 1'd1;
    assign memhint[7668] = 1'd1;
    assign memhint[7669] = 1'd0;
    assign memhint[7670] = 1'd0;
    assign memhint[7671] = 1'd0;
    assign memhint[7672] = 1'd0;
    assign memhint[7673] = 1'd0;
    assign memhint[7674] = 1'd0;
    assign memhint[7675] = 1'd0;
    assign memhint[7676] = 1'd0;
    assign memhint[7677] = 1'd0;
    assign memhint[7678] = 1'd0;
    assign memhint[7679] = 1'd1;
    assign memhint[7680] = 1'd1;
    assign memhint[7681] = 1'd1;
    assign memhint[7682] = 1'd1;
    assign memhint[7683] = 1'd0;
    assign memhint[7684] = 1'd0;
    assign memhint[7685] = 1'd0;
    assign memhint[7686] = 1'd0;
    assign memhint[7687] = 1'd0;
    assign memhint[7688] = 1'd0;
    assign memhint[7689] = 1'd0;
    assign memhint[7690] = 1'd1;
    assign memhint[7691] = 1'd1;
    assign memhint[7692] = 1'd1;
    assign memhint[7693] = 1'd1;
    assign memhint[7694] = 1'd0;
    assign memhint[7695] = 1'd0;
    assign memhint[7696] = 1'd0;
    assign memhint[7697] = 1'd0;
    assign memhint[7698] = 1'd0;
    assign memhint[7699] = 1'd0;
    assign memhint[7700] = 1'd0;
    assign memhint[7701] = 1'd0;
    assign memhint[7702] = 1'd0;
    assign memhint[7703] = 1'd0;
    assign memhint[7704] = 1'd0;
    assign memhint[7705] = 1'd0;
    assign memhint[7706] = 1'd0;
    assign memhint[7707] = 1'd0;
    assign memhint[7708] = 1'd0;
    assign memhint[7709] = 1'd0;
    assign memhint[7710] = 1'd0;
    assign memhint[7711] = 1'd0;
    assign memhint[7712] = 1'd0;
    assign memhint[7713] = 1'd0;
    assign memhint[7714] = 1'd1;
    assign memhint[7715] = 1'd1;
    assign memhint[7716] = 1'd0;
    assign memhint[7717] = 1'd0;
    assign memhint[7718] = 1'd0;
    assign memhint[7719] = 1'd0;
    assign memhint[7720] = 1'd0;
    assign memhint[7721] = 1'd0;
    assign memhint[7722] = 1'd0;
    assign memhint[7723] = 1'd0;
    assign memhint[7724] = 1'd0;
    assign memhint[7725] = 1'd0;
    assign memhint[7726] = 1'd0;
    assign memhint[7727] = 1'd0;
    assign memhint[7728] = 1'd1;
    assign memhint[7729] = 1'd1;
    assign memhint[7730] = 1'd1;
    assign memhint[7731] = 1'd1;
    assign memhint[7732] = 1'd1;
    assign memhint[7733] = 1'd0;
    assign memhint[7734] = 1'd0;
    assign memhint[7735] = 1'd0;
    assign memhint[7736] = 1'd0;
    assign memhint[7737] = 1'd0;
    assign memhint[7738] = 1'd0;
    assign memhint[7739] = 1'd1;
    assign memhint[7740] = 1'd1;
    assign memhint[7741] = 1'd1;
    assign memhint[7742] = 1'd1;
    assign memhint[7743] = 1'd1;
    assign memhint[7744] = 1'd0;
    assign memhint[7745] = 1'd0;
    assign memhint[7746] = 1'd0;
    assign memhint[7747] = 1'd0;
    assign memhint[7748] = 1'd0;
    assign memhint[7749] = 1'd0;
    assign memhint[7750] = 1'd0;
    assign memhint[7751] = 1'd0;
    assign memhint[7752] = 1'd0;
    assign memhint[7753] = 1'd0;
    assign memhint[7754] = 1'd0;
    assign memhint[7755] = 1'd0;
    assign memhint[7756] = 1'd0;
    assign memhint[7757] = 1'd0;
    assign memhint[7758] = 1'd0;
    assign memhint[7759] = 1'd0;
    assign memhint[7760] = 1'd0;
    assign memhint[7761] = 1'd0;
    assign memhint[7762] = 1'd1;
    assign memhint[7763] = 1'd1;
    assign memhint[7764] = 1'd0;
    assign memhint[7765] = 1'd0;
    assign memhint[7766] = 1'd0;
    assign memhint[7767] = 1'd0;
    assign memhint[7768] = 1'd0;
    assign memhint[7769] = 1'd0;
    assign memhint[7770] = 1'd0;
    assign memhint[7771] = 1'd0;
    assign memhint[7772] = 1'd0;
    assign memhint[7773] = 1'd0;
    assign memhint[7774] = 1'd0;
    assign memhint[7775] = 1'd0;
    assign memhint[7776] = 1'd0;
    assign memhint[7777] = 1'd0;
    assign memhint[7778] = 1'd0;
    assign memhint[7779] = 1'd0;
    assign memhint[7780] = 1'd0;
    assign memhint[7781] = 1'd1;
    assign memhint[7782] = 1'd1;
    assign memhint[7783] = 1'd0;
    assign memhint[7784] = 1'd0;
    assign memhint[7785] = 1'd0;
    assign memhint[7786] = 1'd0;
    assign memhint[7787] = 1'd0;
    assign memhint[7788] = 1'd0;
    assign memhint[7789] = 1'd0;
    assign memhint[7790] = 1'd0;
    assign memhint[7791] = 1'd0;
    assign memhint[7792] = 1'd0;
    assign memhint[7793] = 1'd0;
    assign memhint[7794] = 1'd0;
    assign memhint[7795] = 1'd1;
    assign memhint[7796] = 1'd1;
    assign memhint[7797] = 1'd0;
    assign memhint[7798] = 1'd0;
    assign memhint[7799] = 1'd0;
    assign memhint[7800] = 1'd0;
    assign memhint[7801] = 1'd0;
    assign memhint[7802] = 1'd0;
    assign memhint[7803] = 1'd0;
    assign memhint[7804] = 1'd0;
    assign memhint[7805] = 1'd0;
    assign memhint[7806] = 1'd0;
    assign memhint[7807] = 1'd0;
    assign memhint[7808] = 1'd0;
    assign memhint[7809] = 1'd0;
    assign memhint[7810] = 1'd0;
    assign memhint[7811] = 1'd0;
    assign memhint[7812] = 1'd1;
    assign memhint[7813] = 1'd1;
    assign memhint[7814] = 1'd0;
    assign memhint[7815] = 1'd0;
    assign memhint[7816] = 1'd0;
    assign memhint[7817] = 1'd0;
    assign memhint[7818] = 1'd0;
    assign memhint[7819] = 1'd0;
    assign memhint[7820] = 1'd0;
    assign memhint[7821] = 1'd0;
    assign memhint[7822] = 1'd0;
    assign memhint[7823] = 1'd0;
    assign memhint[7824] = 1'd1;
    assign memhint[7825] = 1'd1;
    assign memhint[7826] = 1'd0;
    assign memhint[7827] = 1'd0;
    assign memhint[7828] = 1'd0;
    assign memhint[7829] = 1'd0;
    assign memhint[7830] = 1'd0;
    assign memhint[7831] = 1'd0;
    assign memhint[7832] = 1'd0;
    assign memhint[7833] = 1'd0;
    assign memhint[7834] = 1'd0;
    assign memhint[7835] = 1'd0;
    assign memhint[7836] = 1'd1;
    assign memhint[7837] = 1'd1;
    assign memhint[7838] = 1'd1;
    assign memhint[7839] = 1'd1;
    assign memhint[7840] = 1'd1;
    assign memhint[7841] = 1'd1;
    assign memhint[7842] = 1'd1;
    assign memhint[7843] = 1'd1;
    assign memhint[7844] = 1'd0;
    assign memhint[7845] = 1'd0;
    assign memhint[7846] = 1'd0;
    assign memhint[7847] = 1'd0;
    assign memhint[7848] = 1'd0;
    assign memhint[7849] = 1'd0;
    assign memhint[7850] = 1'd0;
    assign memhint[7851] = 1'd1;
    assign memhint[7852] = 1'd1;
    assign memhint[7853] = 1'd1;
    assign memhint[7854] = 1'd1;
    assign memhint[7855] = 1'd1;
    assign memhint[7856] = 1'd1;
    assign memhint[7857] = 1'd1;
    assign memhint[7858] = 1'd1;
    assign memhint[7859] = 1'd1;
    assign memhint[7860] = 1'd1;
    assign memhint[7861] = 1'd1;
    assign memhint[7862] = 1'd1;
    assign memhint[7863] = 1'd1;
    assign memhint[7864] = 1'd0;
    assign memhint[7865] = 1'd0;
    assign memhint[7866] = 1'd0;
    assign memhint[7867] = 1'd0;
    assign memhint[7868] = 1'd1;
    assign memhint[7869] = 1'd1;
    assign memhint[7870] = 1'd1;
    assign memhint[7871] = 1'd1;
    assign memhint[7872] = 1'd1;
    assign memhint[7873] = 1'd1;
    assign memhint[7874] = 1'd1;
    assign memhint[7875] = 1'd1;
    assign memhint[7876] = 1'd1;
    assign memhint[7877] = 1'd1;
    assign memhint[7878] = 1'd1;
    assign memhint[7879] = 1'd0;
    assign memhint[7880] = 1'd0;
    assign memhint[7881] = 1'd0;
    assign memhint[7882] = 1'd0;
    assign memhint[7883] = 1'd1;
    assign memhint[7884] = 1'd1;
    assign memhint[7885] = 1'd1;
    assign memhint[7886] = 1'd1;
    assign memhint[7887] = 1'd1;
    assign memhint[7888] = 1'd1;
    assign memhint[7889] = 1'd1;
    assign memhint[7890] = 1'd1;
    assign memhint[7891] = 1'd1;
    assign memhint[7892] = 1'd1;
    assign memhint[7893] = 1'd1;
    assign memhint[7894] = 1'd1;
    assign memhint[7895] = 1'd1;
    assign memhint[7896] = 1'd0;
    assign memhint[7897] = 1'd0;
    assign memhint[7898] = 1'd0;
    assign memhint[7899] = 1'd0;
    assign memhint[7900] = 1'd0;
    assign memhint[7901] = 1'd0;
    assign memhint[7902] = 1'd0;
    assign memhint[7903] = 1'd0;
    assign memhint[7904] = 1'd0;
    assign memhint[7905] = 1'd1;
    assign memhint[7906] = 1'd1;
    assign memhint[7907] = 1'd1;
    assign memhint[7908] = 1'd1;
    assign memhint[7909] = 1'd1;
    assign memhint[7910] = 1'd1;
    assign memhint[7911] = 1'd1;
    assign memhint[7912] = 1'd1;
    assign memhint[7913] = 1'd1;
    assign memhint[7914] = 1'd1;
    assign memhint[7915] = 1'd1;
    assign memhint[7916] = 1'd1;
    assign memhint[7917] = 1'd0;
    assign memhint[7918] = 1'd0;
    assign memhint[7919] = 1'd0;
    assign memhint[7920] = 1'd0;
    assign memhint[7921] = 1'd0;
    assign memhint[7922] = 1'd0;
    assign memhint[7923] = 1'd0;
    assign memhint[7924] = 1'd0;
    assign memhint[7925] = 1'd0;
    assign memhint[7926] = 1'd0;
    assign memhint[7927] = 1'd0;
    assign memhint[7928] = 1'd1;
    assign memhint[7929] = 1'd1;
    assign memhint[7930] = 1'd0;
    assign memhint[7931] = 1'd0;
    assign memhint[7932] = 1'd0;
    assign memhint[7933] = 1'd0;
    assign memhint[7934] = 1'd0;
    assign memhint[7935] = 1'd0;
    assign memhint[7936] = 1'd0;
    assign memhint[7937] = 1'd0;
    assign memhint[7938] = 1'd0;
    assign memhint[7939] = 1'd0;
    assign memhint[7940] = 1'd0;
    assign memhint[7941] = 1'd0;
    assign memhint[7942] = 1'd0;
    assign memhint[7943] = 1'd0;
    assign memhint[7944] = 1'd0;
    assign memhint[7945] = 1'd0;
    assign memhint[7946] = 1'd0;
    assign memhint[7947] = 1'd1;
    assign memhint[7948] = 1'd1;
    assign memhint[7949] = 1'd0;
    assign memhint[7950] = 1'd0;
    assign memhint[7951] = 1'd0;
    assign memhint[7952] = 1'd0;
    assign memhint[7953] = 1'd0;
    assign memhint[7954] = 1'd0;
    assign memhint[7955] = 1'd0;
    assign memhint[7956] = 1'd0;
    assign memhint[7957] = 1'd0;
    assign memhint[7958] = 1'd0;
    assign memhint[7959] = 1'd0;
    assign memhint[7960] = 1'd0;
    assign memhint[7961] = 1'd0;
    assign memhint[7962] = 1'd0;
    assign memhint[7963] = 1'd0;
    assign memhint[7964] = 1'd1;
    assign memhint[7965] = 1'd1;
    assign memhint[7966] = 1'd0;
    assign memhint[7967] = 1'd0;
    assign memhint[7968] = 1'd0;
    assign memhint[7969] = 1'd0;
    assign memhint[7970] = 1'd0;
    assign memhint[7971] = 1'd0;
    assign memhint[7972] = 1'd0;
    assign memhint[7973] = 1'd0;
    assign memhint[7974] = 1'd0;
    assign memhint[7975] = 1'd0;
    assign memhint[7976] = 1'd0;
    assign memhint[7977] = 1'd0;
    assign memhint[7978] = 1'd0;
    assign memhint[7979] = 1'd0;
    assign memhint[7980] = 1'd0;
    assign memhint[7981] = 1'd1;
    assign memhint[7982] = 1'd1;
    assign memhint[7983] = 1'd1;
    assign memhint[7984] = 1'd1;
    assign memhint[7985] = 1'd1;
    assign memhint[7986] = 1'd1;
    assign memhint[7987] = 1'd1;
    assign memhint[7988] = 1'd1;
    assign memhint[7989] = 1'd0;
    assign memhint[7990] = 1'd0;
    assign memhint[7991] = 1'd0;
    assign memhint[7992] = 1'd0;
    assign memhint[7993] = 1'd0;
    assign memhint[7994] = 1'd0;
    assign memhint[7995] = 1'd0;
    assign memhint[7996] = 1'd0;
    assign memhint[7997] = 1'd0;
    assign memhint[7998] = 1'd0;
    assign memhint[7999] = 1'd0;
    assign memhint[8000] = 1'd0;
    assign memhint[8001] = 1'd1;
    assign memhint[8002] = 1'd1;
    assign memhint[8003] = 1'd1;
    assign memhint[8004] = 1'd1;
    assign memhint[8005] = 1'd1;
    assign memhint[8006] = 1'd1;
    assign memhint[8007] = 1'd1;
    assign memhint[8008] = 1'd1;
    assign memhint[8009] = 1'd1;
    assign memhint[8010] = 1'd1;
    assign memhint[8011] = 1'd1;
    assign memhint[8012] = 1'd1;
    assign memhint[8013] = 1'd0;
    assign memhint[8014] = 1'd0;
    assign memhint[8015] = 1'd0;
    assign memhint[8016] = 1'd0;
    assign memhint[8017] = 1'd0;
    assign memhint[8018] = 1'd0;
    assign memhint[8019] = 1'd0;
    assign memhint[8020] = 1'd0;
    assign memhint[8021] = 1'd0;
    assign memhint[8022] = 1'd0;
    assign memhint[8023] = 1'd0;
    assign memhint[8024] = 1'd1;
    assign memhint[8025] = 1'd1;
    assign memhint[8026] = 1'd0;
    assign memhint[8027] = 1'd0;
    assign memhint[8028] = 1'd0;
    assign memhint[8029] = 1'd0;
    assign memhint[8030] = 1'd0;
    assign memhint[8031] = 1'd0;
    assign memhint[8032] = 1'd0;
    assign memhint[8033] = 1'd0;
    assign memhint[8034] = 1'd0;
    assign memhint[8035] = 1'd0;
    assign memhint[8036] = 1'd0;
    assign memhint[8037] = 1'd0;
    assign memhint[8038] = 1'd0;
    assign memhint[8039] = 1'd0;
    assign memhint[8040] = 1'd1;
    assign memhint[8041] = 1'd1;
    assign memhint[8042] = 1'd0;
    assign memhint[8043] = 1'd0;
    assign memhint[8044] = 1'd0;
    assign memhint[8045] = 1'd0;
    assign memhint[8046] = 1'd0;
    assign memhint[8047] = 1'd0;
    assign memhint[8048] = 1'd0;
    assign memhint[8049] = 1'd0;
    assign memhint[8050] = 1'd0;
    assign memhint[8051] = 1'd0;
    assign memhint[8052] = 1'd0;
    assign memhint[8053] = 1'd1;
    assign memhint[8054] = 1'd1;
    assign memhint[8055] = 1'd1;
    assign memhint[8056] = 1'd1;
    assign memhint[8057] = 1'd1;
    assign memhint[8058] = 1'd1;
    assign memhint[8059] = 1'd1;
    assign memhint[8060] = 1'd1;
    assign memhint[8061] = 1'd1;
    assign memhint[8062] = 1'd1;
    assign memhint[8063] = 1'd1;
    assign memhint[8064] = 1'd1;
    assign memhint[8065] = 1'd1;
    assign memhint[8066] = 1'd0;
    assign memhint[8067] = 1'd0;
    assign memhint[8068] = 1'd0;
    assign memhint[8069] = 1'd0;
    assign memhint[8070] = 1'd0;
    assign memhint[8071] = 1'd0;
    assign memhint[8072] = 1'd0;
    assign memhint[8073] = 1'd0;
    assign memhint[8074] = 1'd0;
    assign memhint[8075] = 1'd0;
    assign memhint[8076] = 1'd0;
    assign memhint[8077] = 1'd0;
    assign memhint[8078] = 1'd0;
    assign memhint[8079] = 1'd0;
    assign memhint[8080] = 1'd0;
    assign memhint[8081] = 1'd0;
    assign memhint[8082] = 1'd0;
    assign memhint[8083] = 1'd0;
    assign memhint[8084] = 1'd0;
    assign memhint[8085] = 1'd0;
    assign memhint[8086] = 1'd0;
    assign memhint[8087] = 1'd1;
    assign memhint[8088] = 1'd1;
    assign memhint[8089] = 1'd0;
    assign memhint[8090] = 1'd0;
    assign memhint[8091] = 1'd0;
    assign memhint[8092] = 1'd0;
    assign memhint[8093] = 1'd0;
    assign memhint[8094] = 1'd0;
    assign memhint[8095] = 1'd0;
    assign memhint[8096] = 1'd0;
    assign memhint[8097] = 1'd0;
    assign memhint[8098] = 1'd0;
    assign memhint[8099] = 1'd0;
    assign memhint[8100] = 1'd0;
    assign memhint[8101] = 1'd0;
    assign memhint[8102] = 1'd0;
    assign memhint[8103] = 1'd1;
    assign memhint[8104] = 1'd1;
    assign memhint[8105] = 1'd1;
    assign memhint[8106] = 1'd1;
    assign memhint[8107] = 1'd1;
    assign memhint[8108] = 1'd1;
    assign memhint[8109] = 1'd1;
    assign memhint[8110] = 1'd1;
    assign memhint[8111] = 1'd1;
    assign memhint[8112] = 1'd1;
    assign memhint[8113] = 1'd1;
    assign memhint[8114] = 1'd1;
    assign memhint[8115] = 1'd0;
    assign memhint[8116] = 1'd0;
    assign memhint[8117] = 1'd0;
    assign memhint[8118] = 1'd0;
    assign memhint[8119] = 1'd0;
    assign memhint[8120] = 1'd0;
    assign memhint[8121] = 1'd0;
    assign memhint[8122] = 1'd0;
    assign memhint[8123] = 1'd0;
    assign memhint[8124] = 1'd0;
    assign memhint[8125] = 1'd0;
    assign memhint[8126] = 1'd0;
    assign memhint[8127] = 1'd0;
    assign memhint[8128] = 1'd0;
    assign memhint[8129] = 1'd0;
    assign memhint[8130] = 1'd0;
    assign memhint[8131] = 1'd0;
    assign memhint[8132] = 1'd0;
    assign memhint[8133] = 1'd0;
    assign memhint[8134] = 1'd0;
    assign memhint[8135] = 1'd1;
    assign memhint[8136] = 1'd1;
    assign memhint[8137] = 1'd0;
    assign memhint[8138] = 1'd0;
    assign memhint[8139] = 1'd0;
    assign memhint[8140] = 1'd0;
    assign memhint[8141] = 1'd0;
    assign memhint[8142] = 1'd0;
    assign memhint[8143] = 1'd0;
    assign memhint[8144] = 1'd0;
    assign memhint[8145] = 1'd0;
    assign memhint[8146] = 1'd0;
    assign memhint[8147] = 1'd0;
    assign memhint[8148] = 1'd0;
    assign memhint[8149] = 1'd0;
    assign memhint[8150] = 1'd0;
    assign memhint[8151] = 1'd0;
    assign memhint[8152] = 1'd0;
    assign memhint[8153] = 1'd0;
    assign memhint[8154] = 1'd1;
    assign memhint[8155] = 1'd1;
    assign memhint[8156] = 1'd1;
    assign memhint[8157] = 1'd1;
    assign memhint[8158] = 1'd1;
    assign memhint[8159] = 1'd1;
    assign memhint[8160] = 1'd1;
    assign memhint[8161] = 1'd1;
    assign memhint[8162] = 1'd1;
    assign memhint[8163] = 1'd1;
    assign memhint[8164] = 1'd1;
    assign memhint[8165] = 1'd0;
    assign memhint[8166] = 1'd0;
    assign memhint[8167] = 1'd0;
    assign memhint[8168] = 1'd1;
    assign memhint[8169] = 1'd1;
    assign memhint[8170] = 1'd0;
    assign memhint[8171] = 1'd0;
    assign memhint[8172] = 1'd0;
    assign memhint[8173] = 1'd0;
    assign memhint[8174] = 1'd0;
    assign memhint[8175] = 1'd0;
    assign memhint[8176] = 1'd0;
    assign memhint[8177] = 1'd0;
    assign memhint[8178] = 1'd0;
    assign memhint[8179] = 1'd0;
    assign memhint[8180] = 1'd0;
    assign memhint[8181] = 1'd0;
    assign memhint[8182] = 1'd0;
    assign memhint[8183] = 1'd0;
    assign memhint[8184] = 1'd0;
    assign memhint[8185] = 1'd1;
    assign memhint[8186] = 1'd1;
    assign memhint[8187] = 1'd0;
    assign memhint[8188] = 1'd0;
    assign memhint[8189] = 1'd0;
    assign memhint[8190] = 1'd0;
    assign memhint[8191] = 1'd0;
    assign memhint[8192] = 1'd0;
    assign memhint[8193] = 1'd0;
    assign memhint[8194] = 1'd0;
    assign memhint[8195] = 1'd0;
    assign memhint[8196] = 1'd0;
    assign memhint[8197] = 1'd1;
    assign memhint[8198] = 1'd1;
    assign memhint[8199] = 1'd0;
    assign memhint[8200] = 1'd0;
    assign memhint[8201] = 1'd0;
    assign memhint[8202] = 1'd0;
    assign memhint[8203] = 1'd0;
    assign memhint[8204] = 1'd0;
    assign memhint[8205] = 1'd0;
    assign memhint[8206] = 1'd0;
    assign memhint[8207] = 1'd0;
    assign memhint[8208] = 1'd0;
    assign memhint[8209] = 1'd0;
    assign memhint[8210] = 1'd1;
    assign memhint[8211] = 1'd1;
    assign memhint[8212] = 1'd1;
    assign memhint[8213] = 1'd1;
    assign memhint[8214] = 1'd1;
    assign memhint[8215] = 1'd0;
    assign memhint[8216] = 1'd0;
    assign memhint[8217] = 1'd0;
    assign memhint[8218] = 1'd0;
    assign memhint[8219] = 1'd0;
    assign memhint[8220] = 1'd0;
    assign memhint[8221] = 1'd0;
    assign memhint[8222] = 1'd0;
    assign memhint[8223] = 1'd0;
    assign memhint[8224] = 1'd1;
    assign memhint[8225] = 1'd1;
    assign memhint[8226] = 1'd1;
    assign memhint[8227] = 1'd1;
    assign memhint[8228] = 1'd1;
    assign memhint[8229] = 1'd1;
    assign memhint[8230] = 1'd1;
    assign memhint[8231] = 1'd1;
    assign memhint[8232] = 1'd1;
    assign memhint[8233] = 1'd1;
    assign memhint[8234] = 1'd1;
    assign memhint[8235] = 1'd1;
    assign memhint[8236] = 1'd1;
    assign memhint[8237] = 1'd0;
    assign memhint[8238] = 1'd0;
    assign memhint[8239] = 1'd0;
    assign memhint[8240] = 1'd0;
    assign memhint[8241] = 1'd1;
    assign memhint[8242] = 1'd1;
    assign memhint[8243] = 1'd1;
    assign memhint[8244] = 1'd1;
    assign memhint[8245] = 1'd1;
    assign memhint[8246] = 1'd1;
    assign memhint[8247] = 1'd1;
    assign memhint[8248] = 1'd1;
    assign memhint[8249] = 1'd1;
    assign memhint[8250] = 1'd1;
    assign memhint[8251] = 1'd1;
    assign memhint[8252] = 1'd0;
    assign memhint[8253] = 1'd0;
    assign memhint[8254] = 1'd0;
    assign memhint[8255] = 1'd0;
    assign memhint[8256] = 1'd1;
    assign memhint[8257] = 1'd1;
    assign memhint[8258] = 1'd1;
    assign memhint[8259] = 1'd1;
    assign memhint[8260] = 1'd1;
    assign memhint[8261] = 1'd1;
    assign memhint[8262] = 1'd1;
    assign memhint[8263] = 1'd1;
    assign memhint[8264] = 1'd1;
    assign memhint[8265] = 1'd1;
    assign memhint[8266] = 1'd1;
    assign memhint[8267] = 1'd1;
    assign memhint[8268] = 1'd1;
    assign memhint[8269] = 1'd0;
    assign memhint[8270] = 1'd0;
    assign memhint[8271] = 1'd0;
    assign memhint[8272] = 1'd0;
    assign memhint[8273] = 1'd0;
    assign memhint[8274] = 1'd0;
    assign memhint[8275] = 1'd0;
    assign memhint[8276] = 1'd0;
    assign memhint[8277] = 1'd0;
    assign memhint[8278] = 1'd0;
    assign memhint[8279] = 1'd0;
    assign memhint[8280] = 1'd1;
    assign memhint[8281] = 1'd1;
    assign memhint[8282] = 1'd1;
    assign memhint[8283] = 1'd1;
    assign memhint[8284] = 1'd1;
    assign memhint[8285] = 1'd1;
    assign memhint[8286] = 1'd1;
    assign memhint[8287] = 1'd1;
    assign memhint[8288] = 1'd0;
    assign memhint[8289] = 1'd0;
    assign memhint[8290] = 1'd0;
    assign memhint[8291] = 1'd0;
    assign memhint[8292] = 1'd0;
    assign memhint[8293] = 1'd0;
    assign memhint[8294] = 1'd0;
    assign memhint[8295] = 1'd0;
    assign memhint[8296] = 1'd0;
    assign memhint[8297] = 1'd0;
    assign memhint[8298] = 1'd0;
    assign memhint[8299] = 1'd0;
    assign memhint[8300] = 1'd0;
    assign memhint[8301] = 1'd1;
    assign memhint[8302] = 1'd1;
    assign memhint[8303] = 1'd0;
    assign memhint[8304] = 1'd0;
    assign memhint[8305] = 1'd0;
    assign memhint[8306] = 1'd0;
    assign memhint[8307] = 1'd0;
    assign memhint[8308] = 1'd0;
    assign memhint[8309] = 1'd0;
    assign memhint[8310] = 1'd0;
    assign memhint[8311] = 1'd0;
    assign memhint[8312] = 1'd0;
    assign memhint[8313] = 1'd0;
    assign memhint[8314] = 1'd0;
    assign memhint[8315] = 1'd0;
    assign memhint[8316] = 1'd0;
    assign memhint[8317] = 1'd0;
    assign memhint[8318] = 1'd0;
    assign memhint[8319] = 1'd1;
    assign memhint[8320] = 1'd1;
    assign memhint[8321] = 1'd0;
    assign memhint[8322] = 1'd0;
    assign memhint[8323] = 1'd0;
    assign memhint[8324] = 1'd0;
    assign memhint[8325] = 1'd0;
    assign memhint[8326] = 1'd0;
    assign memhint[8327] = 1'd0;
    assign memhint[8328] = 1'd0;
    assign memhint[8329] = 1'd0;
    assign memhint[8330] = 1'd0;
    assign memhint[8331] = 1'd0;
    assign memhint[8332] = 1'd0;
    assign memhint[8333] = 1'd0;
    assign memhint[8334] = 1'd0;
    assign memhint[8335] = 1'd0;
    assign memhint[8336] = 1'd0;
    assign memhint[8337] = 1'd0;
    assign memhint[8338] = 1'd1;
    assign memhint[8339] = 1'd1;
    assign memhint[8340] = 1'd0;
    assign memhint[8341] = 1'd0;
    assign memhint[8342] = 1'd0;
    assign memhint[8343] = 1'd0;
    assign memhint[8344] = 1'd0;
    assign memhint[8345] = 1'd0;
    assign memhint[8346] = 1'd0;
    assign memhint[8347] = 1'd0;
    assign memhint[8348] = 1'd0;
    assign memhint[8349] = 1'd0;
    assign memhint[8350] = 1'd0;
    assign memhint[8351] = 1'd0;
    assign memhint[8352] = 1'd0;
    assign memhint[8353] = 1'd0;
    assign memhint[8354] = 1'd0;
    assign memhint[8355] = 1'd1;
    assign memhint[8356] = 1'd1;
    assign memhint[8357] = 1'd1;
    assign memhint[8358] = 1'd1;
    assign memhint[8359] = 1'd1;
    assign memhint[8360] = 1'd0;
    assign memhint[8361] = 1'd0;
    assign memhint[8362] = 1'd0;
    assign memhint[8363] = 1'd0;
    assign memhint[8364] = 1'd0;
    assign memhint[8365] = 1'd0;
    assign memhint[8366] = 1'd0;
    assign memhint[8367] = 1'd0;
    assign memhint[8368] = 1'd0;
    assign memhint[8369] = 1'd0;
    assign memhint[8370] = 1'd0;
    assign memhint[8371] = 1'd0;
    assign memhint[8372] = 1'd0;
    assign memhint[8373] = 1'd0;
    assign memhint[8374] = 1'd0;
    assign memhint[8375] = 1'd0;
    assign memhint[8376] = 1'd1;
    assign memhint[8377] = 1'd1;
    assign memhint[8378] = 1'd1;
    assign memhint[8379] = 1'd1;
    assign memhint[8380] = 1'd1;
    assign memhint[8381] = 1'd1;
    assign memhint[8382] = 1'd1;
    assign memhint[8383] = 1'd1;
    assign memhint[8384] = 1'd0;
    assign memhint[8385] = 1'd0;
    assign memhint[8386] = 1'd0;
    assign memhint[8387] = 1'd0;
    assign memhint[8388] = 1'd0;
    assign memhint[8389] = 1'd0;
    assign memhint[8390] = 1'd0;
    assign memhint[8391] = 1'd0;
    assign memhint[8392] = 1'd0;
    assign memhint[8393] = 1'd0;
    assign memhint[8394] = 1'd0;
    assign memhint[8395] = 1'd0;
    assign memhint[8396] = 1'd0;
    assign memhint[8397] = 1'd1;
    assign memhint[8398] = 1'd1;
    assign memhint[8399] = 1'd0;
    assign memhint[8400] = 1'd0;
    assign memhint[8401] = 1'd0;
    assign memhint[8402] = 1'd0;
    assign memhint[8403] = 1'd0;
    assign memhint[8404] = 1'd0;
    assign memhint[8405] = 1'd0;
    assign memhint[8406] = 1'd0;
    assign memhint[8407] = 1'd0;
    assign memhint[8408] = 1'd0;
    assign memhint[8409] = 1'd0;
    assign memhint[8410] = 1'd0;
    assign memhint[8411] = 1'd0;
    assign memhint[8412] = 1'd0;
    assign memhint[8413] = 1'd0;
    assign memhint[8414] = 1'd1;
    assign memhint[8415] = 1'd0;
    assign memhint[8416] = 1'd0;
    assign memhint[8417] = 1'd0;
    assign memhint[8418] = 1'd0;
    assign memhint[8419] = 1'd0;
    assign memhint[8420] = 1'd0;
    assign memhint[8421] = 1'd0;
    assign memhint[8422] = 1'd0;
    assign memhint[8423] = 1'd0;
    assign memhint[8424] = 1'd0;
    assign memhint[8425] = 1'd0;
    assign memhint[8426] = 1'd0;
    assign memhint[8427] = 1'd0;
    assign memhint[8428] = 1'd0;
    assign memhint[8429] = 1'd1;
    assign memhint[8430] = 1'd1;
    assign memhint[8431] = 1'd1;
    assign memhint[8432] = 1'd1;
    assign memhint[8433] = 1'd1;
    assign memhint[8434] = 1'd1;
    assign memhint[8435] = 1'd1;
    assign memhint[8436] = 1'd1;
    assign memhint[8437] = 1'd0;
    assign memhint[8438] = 1'd0;
    assign memhint[8439] = 1'd0;
    assign memhint[8440] = 1'd0;
    assign memhint[8441] = 1'd0;
    assign memhint[8442] = 1'd0;
    assign memhint[8443] = 1'd0;
    assign memhint[8444] = 1'd0;
    assign memhint[8445] = 1'd0;
    assign memhint[8446] = 1'd0;
    assign memhint[8447] = 1'd0;
    assign memhint[8448] = 1'd0;
    assign memhint[8449] = 1'd0;
    assign memhint[8450] = 1'd0;
    assign memhint[8451] = 1'd0;
    assign memhint[8452] = 1'd0;
    assign memhint[8453] = 1'd0;
    assign memhint[8454] = 1'd0;
    assign memhint[8455] = 1'd0;
    assign memhint[8456] = 1'd0;
    assign memhint[8457] = 1'd0;
    assign memhint[8458] = 1'd0;
    assign memhint[8459] = 1'd0;
    assign memhint[8460] = 1'd1;
    assign memhint[8461] = 1'd1;
    assign memhint[8462] = 1'd0;
    assign memhint[8463] = 1'd0;
    assign memhint[8464] = 1'd0;
    assign memhint[8465] = 1'd0;
    assign memhint[8466] = 1'd0;
    assign memhint[8467] = 1'd0;
    assign memhint[8468] = 1'd0;
    assign memhint[8469] = 1'd0;
    assign memhint[8470] = 1'd0;
    assign memhint[8471] = 1'd0;
    assign memhint[8472] = 1'd0;
    assign memhint[8473] = 1'd0;
    assign memhint[8474] = 1'd0;
    assign memhint[8475] = 1'd0;
    assign memhint[8476] = 1'd0;
    assign memhint[8477] = 1'd0;
    assign memhint[8478] = 1'd1;
    assign memhint[8479] = 1'd1;
    assign memhint[8480] = 1'd1;
    assign memhint[8481] = 1'd1;
    assign memhint[8482] = 1'd1;
    assign memhint[8483] = 1'd1;
    assign memhint[8484] = 1'd1;
    assign memhint[8485] = 1'd1;
    assign memhint[8486] = 1'd0;
    assign memhint[8487] = 1'd0;
    assign memhint[8488] = 1'd0;
    assign memhint[8489] = 1'd0;
    assign memhint[8490] = 1'd0;
    assign memhint[8491] = 1'd0;
    assign memhint[8492] = 1'd0;
    assign memhint[8493] = 1'd0;
    assign memhint[8494] = 1'd0;
    assign memhint[8495] = 1'd0;
    assign memhint[8496] = 1'd0;
    assign memhint[8497] = 1'd0;
    assign memhint[8498] = 1'd0;
    assign memhint[8499] = 1'd0;
    assign memhint[8500] = 1'd0;
    assign memhint[8501] = 1'd0;
    assign memhint[8502] = 1'd0;
    assign memhint[8503] = 1'd0;
    assign memhint[8504] = 1'd0;
    assign memhint[8505] = 1'd0;
    assign memhint[8506] = 1'd0;
    assign memhint[8507] = 1'd0;
    assign memhint[8508] = 1'd1;
    assign memhint[8509] = 1'd1;
    assign memhint[8510] = 1'd0;
    assign memhint[8511] = 1'd0;
    assign memhint[8512] = 1'd0;
    assign memhint[8513] = 1'd0;
    assign memhint[8514] = 1'd0;
    assign memhint[8515] = 1'd0;
    assign memhint[8516] = 1'd0;
    assign memhint[8517] = 1'd0;
    assign memhint[8518] = 1'd0;
    assign memhint[8519] = 1'd0;
    assign memhint[8520] = 1'd0;
    assign memhint[8521] = 1'd0;
    assign memhint[8522] = 1'd0;
    assign memhint[8523] = 1'd0;
    assign memhint[8524] = 1'd0;
    assign memhint[8525] = 1'd0;
    assign memhint[8526] = 1'd0;
    assign memhint[8527] = 1'd1;
    assign memhint[8528] = 1'd1;
    assign memhint[8529] = 1'd1;
    assign memhint[8530] = 1'd1;
    assign memhint[8531] = 1'd1;
    assign memhint[8532] = 1'd1;
    assign memhint[8533] = 1'd1;
    assign memhint[8534] = 1'd1;
    assign memhint[8535] = 1'd1;
    assign memhint[8536] = 1'd1;
    assign memhint[8537] = 1'd1;
    assign memhint[8538] = 1'd0;
    assign memhint[8539] = 1'd0;
    assign memhint[8540] = 1'd1;
    assign memhint[8541] = 1'd1;
    assign memhint[8542] = 1'd0;
    assign memhint[8543] = 1'd0;
    assign memhint[8544] = 1'd0;
    assign memhint[8545] = 1'd0;
    assign memhint[8546] = 1'd0;
    assign memhint[8547] = 1'd0;
    assign memhint[8548] = 1'd0;
    assign memhint[8549] = 1'd0;
    assign memhint[8550] = 1'd0;
    assign memhint[8551] = 1'd0;
    assign memhint[8552] = 1'd0;
    assign memhint[8553] = 1'd0;
    assign memhint[8554] = 1'd0;
    assign memhint[8555] = 1'd0;
    assign memhint[8556] = 1'd0;
    assign memhint[8557] = 1'd0;
    assign memhint[8558] = 1'd0;
    assign memhint[8559] = 1'd1;
    assign memhint[8560] = 1'd1;
    assign memhint[8561] = 1'd0;
    assign memhint[8562] = 1'd0;
    assign memhint[8563] = 1'd0;
    assign memhint[8564] = 1'd0;
    assign memhint[8565] = 1'd0;
    assign memhint[8566] = 1'd0;
    assign memhint[8567] = 1'd0;
    assign memhint[8568] = 1'd0;
    assign memhint[8569] = 1'd0;
    assign memhint[8570] = 1'd1;
    assign memhint[8571] = 1'd1;
    assign memhint[8572] = 1'd0;
    assign memhint[8573] = 1'd0;
    assign memhint[8574] = 1'd0;
    assign memhint[8575] = 1'd0;
    assign memhint[8576] = 1'd0;
    assign memhint[8577] = 1'd0;
    assign memhint[8578] = 1'd0;

endmodule
