//	How to use:	
//	1. Edit the songs on the Enter Song sheet.	
// 	2. Select this whole worksheet, copy it, and paste it into a new file.	
//	3. Save the file as song_rom.v.	

module pulse1_rom (
    input clk,						
	output reg [25:0] dout,						
	input [11:0] addr		
    );
        
    wire [25:0] memory [4095:0];  			
	always @(posedge clk)						
		dout = memory[addr];					

    parameter s1 = 526;
    parameter s2 = s1 + 291;
    parameter s3 = s2 + 81;

    assign memory[0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[1  ] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[2  ] = {7'd49 , 8'd96 , 7'd85 , 2'd1, 2'd0};   //note: 5A
    assign memory[3  ] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[4  ] = {7'd47 , 8'd96 , 7'd84 , 2'd1, 2'd0};   //note: 5G
    assign memory[5  ] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[6  ] = {7'd49 , 8'd96 , 7'd84 , 2'd1, 2'd0};   //note: 5A
    assign memory[7  ] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[8  ] = {7'd47 , 8'd96 , 7'd83 , 2'd1, 2'd0};   //note: 5G
    assign memory[9  ] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[10 ] = {7'd49 , 8'd96 , 7'd83 , 2'd1, 2'd0};   //note: 5A
    assign memory[11 ] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[12 ] = {7'd47 , 8'd96 , 7'd83 , 2'd1, 2'd0};   //note: 5G
    assign memory[13 ] = {7'd49 , 8'd48 , 7'd83 , 2'd1, 2'd0};   //note: 5A
    assign memory[14 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[15 ] = {7'd49 , 8'd48 , 7'd83 , 2'd1, 2'd0};   //note: 5A
    assign memory[16 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[17 ] = {7'd47 , 8'd48 , 7'd83 , 2'd1, 2'd0};   //note: 5G
    assign memory[18 ] = {7'd49 , 8'd48 , 7'd83 , 2'd1, 2'd0};   //note: 5A
    assign memory[19 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[20 ] = {7'd50 , 8'd96 , 7'd83 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[21 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[22 ] = {7'd49 , 8'd48 , 7'd84 , 2'd1, 2'd0};   //note: 5A
    assign memory[23 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[24 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[25 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[26 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[27 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[28 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[29 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[30 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[31 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[32 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[33 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[34 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[35 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[36 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[37 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[38 ] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[39 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[40 ] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[41 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[42 ] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[43 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[44 ] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[45 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[46 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[47 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[48 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[49 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[50 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[51 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[52 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[53 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[54 ] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[55 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[56 ] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[57 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[58 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[59 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[60 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[61 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[62 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[63 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[64 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[65 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[66 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[67 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[68 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[69 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[70 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[71 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[72 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[73 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[74 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[75 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[76 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[77 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[78 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[79 ] = {7'd48 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G#Ab
    assign memory[80 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[81 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[82 ] = {7'd46 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F#Gb
    assign memory[83 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[84 ] = {7'd47 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[85 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[86 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[87 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[88 ] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[89 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[90 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[91 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[92 ] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[93 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[94 ] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[95 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[96 ] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[97 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[98 ] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[99 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[100] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[101] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[102] = {7'd54 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6D
    assign memory[103] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[104] = {7'd54 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6D
    assign memory[105] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[106] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[107] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[108] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[109] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[110] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[111] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[112] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[113] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[114] = {7'd55 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[115] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[116] = {7'd55 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[117] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[118] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[119] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[120] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[121] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[122] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[123] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[124] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[125] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[126] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[127] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[128] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[129] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[130] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[131] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[132] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[133] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[134] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[135] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[136] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[137] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[138] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[139] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[140] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[141] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[142] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[143] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[144] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[145] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[146] = {7'd44 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5E
    assign memory[147] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[148] = {7'd44 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5E
    assign memory[149] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[150] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[151] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[152] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[153] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[154] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[155] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[156] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[157] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[158] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[159] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[160] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[161] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[162] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[163] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[164] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[165] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[166] = {7'd54 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6D
    assign memory[167] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[168] = {7'd54 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6D
    assign memory[169] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[170] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[171] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[172] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[173] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[174] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[175] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[176] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[177] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[178] = {7'd55 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[179] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[180] = {7'd55 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[181] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[182] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[183] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[184] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[185] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[186] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[187] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[188] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[189] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[190] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[191] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[192] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[193] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[194] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[195] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[196] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[197] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[198] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[199] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[200] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[201] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[202] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[203] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[204] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[205] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[206] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[207] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[208] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[209] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[210] = {7'd56 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6E
    assign memory[211] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[212] = {7'd56 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6E
    assign memory[213] = {7'd45 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[214] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[215] = {7'd45 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[216] = {7'd47 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[217] = {7'd49 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[218] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[219] = {7'd47 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[220] = {7'd52 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[221] = {7'd45 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[222] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[223] = {7'd45 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[224] = {7'd44 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5E
    assign memory[225] = {7'd49 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[226] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[227] = {7'd47 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[228] = {7'd52 , 8'd192, 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[229] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[230] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[231] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[232] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[233] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[234] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[235] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[236] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[237] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[238] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[239] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[240] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[241] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[242] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[243] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[244] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[245] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[246] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[247] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[248] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[249] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[250] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[251] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[252] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[253] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[254] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[255] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[256] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[257] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[258] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[259] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[260] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[261] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[262] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[263] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[264] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[265] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[266] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[267] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[268] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[269] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[270] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[271] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[272] = {7'd45 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F
    assign memory[273] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[274] = {7'd44 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5E
    assign memory[275] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[276] = {7'd44 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5E
    assign memory[277] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[278] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[279] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[280] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[281] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[282] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[283] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[284] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[285] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[286] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[287] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[288] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[289] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[290] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[291] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[292] = {7'd52 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 6C
    assign memory[293] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[294] = {7'd49 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[295] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[296] = {7'd47 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[297] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[298] = {7'd49 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[299] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[300] = {7'd47 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[301] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[302] = {7'd49 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[303] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[304] = {7'd47 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[305] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[306] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[307] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[308] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[309] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[310] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[311] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[312] = {7'd50 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[313] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[314] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[315] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[316] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[317] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[318] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[319] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[320] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[321] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[322] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[323] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[324] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[325] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[326] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[327] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[328] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[329] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[330] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[331] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[332] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[333] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[334] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[335] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[336] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[337] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[338] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[339] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[340] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[341] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[342] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[343] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[344] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[345] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[346] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[347] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[348] = {7'd50 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[349] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[350] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[351] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[352] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[353] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[354] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[355] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[356] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[357] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[358] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[359] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[360] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[361] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[362] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[363] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[364] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[365] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[366] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[367] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[368] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[369] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[370] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[371] = {7'd48 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G#Ab
    assign memory[372] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[373] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[374] = {7'd46 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5F#Gb
    assign memory[375] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[376] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[377] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[378] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[379] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[380] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[381] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[382] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[383] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[384] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[385] = {7'd54 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D
    assign memory[386] = {7'd54 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D
    assign memory[387] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[388] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[389] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[390] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[391] = {7'd55 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[392] = {7'd55 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[393] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[394] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[395] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[396] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[397] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[398] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[399] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[400] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[401] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[402] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[403] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[404] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[405] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[406] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[407] = {7'd44 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5E
    assign memory[408] = {7'd44 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5E
    assign memory[409] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[410] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[411] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[412] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[413] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[414] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[415] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[416] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[417] = {7'd54 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D
    assign memory[418] = {7'd54 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D
    assign memory[419] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[420] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[421] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[422] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[423] = {7'd55 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[424] = {7'd55 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[425] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[426] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[427] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[428] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[429] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[430] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[431] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[432] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[433] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[434] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[435] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[436] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[437] = {7'd52 , 8'd72 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[438] = {7'd52 , 8'd72 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[439] = {7'd52 , 8'd48 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[440] = {7'd56 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6E
    assign memory[441] = {7'd56 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6E
    assign memory[442] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[443] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[444] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[445] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[446] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[447] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[448] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[449] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[450] = {7'd54 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D
    assign memory[451] = {7'd54 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D
    assign memory[452] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[453] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[454] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[455] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[456] = {7'd55 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[457] = {7'd55 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[458] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[459] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[460] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[461] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[462] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[463] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[464] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[465] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[466] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[467] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[468] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[469] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[470] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[471] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[472] = {7'd44 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5E
    assign memory[473] = {7'd44 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5E
    assign memory[474] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[475] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[476] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[477] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[478] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[479] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[480] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[481] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[482] = {7'd54 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D
    assign memory[483] = {7'd54 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D
    assign memory[484] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[485] = {7'd50 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A#Bb
    assign memory[486] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[487] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[488] = {7'd55 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[489] = {7'd55 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6D#Eb
    assign memory[490] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[491] = {7'd49 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5A
    assign memory[492] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[493] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[494] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[495] = {7'd52 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[496] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[497] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[498] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[499] = {7'd45 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5F
    assign memory[500] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[501] = {7'd47 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 5G
    assign memory[502] = {7'd52 , 8'd72 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[503] = {7'd52 , 8'd72 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[504] = {7'd52 , 8'd48 , 7'd106, 2'd1, 2'd0};   //note: 6C
    assign memory[505] = {7'd56 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6E
    assign memory[506] = {7'd56 , 8'd96 , 7'd106, 2'd1, 2'd0};   //note: 6E
    assign memory[507] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[508] = {7'd49 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[509] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[510] = {7'd47 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[511] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[512] = {7'd49 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[513] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[514] = {7'd47 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[515] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[516] = {7'd49 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[517] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[518] = {7'd47 , 8'd96 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[519] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[520] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[521] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[522] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[523] = {7'd47 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5G
    assign memory[524] = {7'd49 , 8'd48 , 7'd96 , 2'd1, 2'd0};   //note: 5A
    assign memory[525] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s1+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s1+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+13 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+14 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+15 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+16 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+17 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+18 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+19 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+20 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+21 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+22 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+23 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+24 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+25 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+26 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+27 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+28 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+29 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+30 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+31 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+32 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+33 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+34 ] = {7'd34 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+35 ] = {7'd36 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+36 ] = {7'd34 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+37 ] = {7'd36 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+38 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+39 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+40 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+41 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+42 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+43 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+44 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+45 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+46 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+47 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+48 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+49 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+50 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+51 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+52 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+53 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+54 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+55 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+56 ] = {7'd36 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+57 ] = {7'd34 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+58 ] = {7'd36 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+59 ] = {7'd34 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+60 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+61 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+62 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+63 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+64 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+65 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+66 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+67 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+68 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+69 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+70 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+71 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+72 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+73 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+74 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+75 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+76 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+77 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+78 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+79 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+80 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+81 ] = {7'd34 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+82 ] = {7'd36 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+83 ] = {7'd34 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+84 ] = {7'd36 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+85 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+86 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+87 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+88 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+89 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+90 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+91 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+92 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+93 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+94 ] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+95 ] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+96 ] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+97 ] = {7'd19 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+98 ] = {7'd19 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3D#Eb
    assign memory[s1+99 ] = {7'd26 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s1+100] = {7'd31 , 8'd48 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+101] = {7'd29 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+102] = {7'd31 , 8'd24 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+103] = {7'd36 , 8'd32 , 7'd123, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+104] = {7'd34 , 8'd32 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+105] = {7'd36 , 8'd32 , 7'd123, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+106] = {7'd34 , 8'd32 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+107] = {7'd31 , 8'd32 , 7'd123, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+108] = {7'd34 , 8'd32 , 7'd123, 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+109] = {7'd31 , 8'd96 , 7'd46 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+110] = {7'd0  , 8'd240, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+111] = {7'd31 , 8'd24 , 7'd42 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+112] = {7'd31 , 8'd24 , 7'd42 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+113] = {7'd31 , 8'd96 , 7'd41 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+114] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+115] = {7'd0  , 8'd33 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+116] = {7'd31 , 8'd96 , 7'd46 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+117] = {7'd0  , 8'd240, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+118] = {7'd31 , 8'd24 , 7'd46 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+119] = {7'd31 , 8'd24 , 7'd46 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+120] = {7'd31 , 8'd96 , 7'd48 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+121] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+122] = {7'd0  , 8'd33 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+123] = {7'd31 , 8'd96 , 7'd48 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+124] = {7'd0  , 8'd240, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+125] = {7'd31 , 8'd24 , 7'd48 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+126] = {7'd31 , 8'd24 , 7'd48 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+127] = {7'd31 , 8'd96 , 7'd49 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+128] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+129] = {7'd0  , 8'd33 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+130] = {7'd31 , 8'd96 , 7'd48 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+131] = {7'd0  , 8'd240, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+132] = {7'd31 , 8'd24 , 7'd48 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+133] = {7'd31 , 8'd24 , 7'd47 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+134] = {7'd31 , 8'd96 , 7'd47 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+135] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+136] = {7'd36 , 8'd32 , 7'd47 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+137] = {7'd34 , 8'd32 , 7'd42 , 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+138] = {7'd36 , 8'd32 , 7'd42 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s1+139] = {7'd34 , 8'd32 , 7'd41 , 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+140] = {7'd31 , 8'd32 , 7'd41 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+141] = {7'd34 , 8'd32 , 7'd41 , 2'd0, 2'd0};   //note: 4F#Gb
    assign memory[s1+142] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+143] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+144] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+145] = {7'd31 , 8'd3  , 7'd100, 2'd0, 2'd0};
    assign memory[s1+146] = {7'd27 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+147] = {7'd27 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+148] = {7'd29 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+149] = {7'd30 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+150] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+151] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+152] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+153] = {7'd31 , 8'd3  , 7'd100, 2'd0, 2'd0};
    assign memory[s1+154] = {7'd27 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+155] = {7'd27 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+156] = {7'd29 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+157] = {7'd30 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+158] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+159] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+160] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+161] = {7'd31 , 8'd3  , 7'd100, 2'd0, 2'd0};
    assign memory[s1+162] = {7'd27 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+163] = {7'd27 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+164] = {7'd29 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+165] = {7'd30 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+166] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+167] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+168] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+169] = {7'd31 , 8'd3  , 7'd100, 2'd0, 2'd0};
    assign memory[s1+170] = {7'd27 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+171] = {7'd27 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+172] = {7'd29 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+173] = {7'd30 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+174] = {7'd27 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+175] = {7'd27 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+176] = {7'd29 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+177] = {7'd29 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+178] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+179] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+180] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+181] = {7'd31 , 8'd3  , 7'd100, 2'd0, 2'd0};
    assign memory[s1+182] = {7'd27 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+183] = {7'd27 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+184] = {7'd29 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+185] = {7'd29 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+186] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+187] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+188] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+189] = {7'd31 , 8'd3  , 7'd100, 2'd0, 2'd0};
    assign memory[s1+190] = {7'd27 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+191] = {7'd27 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+192] = {7'd29 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+193] = {7'd29 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+194] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+195] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+196] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};
    assign memory[s1+197] = {7'd31 , 8'd3  , 7'd100, 2'd0, 2'd0};
    assign memory[s1+198] = {7'd27 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+199] = {7'd27 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+200] = {7'd29 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+201] = {7'd29 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s1+202] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+203] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+204] = {7'd0  , 8'd66 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+205] = {7'd31 , 8'd192, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+206] = {7'd27 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+207] = {7'd27 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+208] = {7'd29 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+209] = {7'd29 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+210] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+211] = {7'd31 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+212] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+213] = {7'd31 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+214] = {7'd27 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+215] = {7'd27 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+216] = {7'd29 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+217] = {7'd29 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+218] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+219] = {7'd31 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+220] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+221] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+222] = {7'd28 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+223] = {7'd28 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+224] = {7'd30 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+225] = {7'd30 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+226] = {7'd32 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+227] = {7'd32 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+228] = {7'd32 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+229] = {7'd32 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+230] = {7'd28 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4C
    assign memory[s1+231] = {7'd28 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+232] = {7'd30 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D
    assign memory[s1+233] = {7'd30 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+234] = {7'd32 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+235] = {7'd32 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+236] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+237] = {7'd32 , 8'd192, 7'd112, 2'd0, 2'd0};   //note: 4E
    assign memory[s1+238] = {7'd32 , 8'd72 , 7'd98 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+239] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+240] = {7'd32 , 8'd57 , 7'd93 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+241] = {7'd0  , 8'd7  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+242] = {7'd32 , 8'd44 , 7'd88 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+243] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+244] = {7'd32 , 8'd72 , 7'd85 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+245] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+246] = {7'd32 , 8'd57 , 7'd80 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+247] = {7'd0  , 8'd7  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+248] = {7'd32 , 8'd44 , 7'd76 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+249] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+250] = {7'd32 , 8'd72 , 7'd73 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+251] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+252] = {7'd32 , 8'd57 , 7'd68 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+253] = {7'd0  , 8'd7  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+254] = {7'd32 , 8'd44 , 7'd62 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+255] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+256] = {7'd32 , 8'd72 , 7'd55 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+257] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+258] = {7'd32 , 8'd57 , 7'd52 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+259] = {7'd0  , 8'd7  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+260] = {7'd32 , 8'd44 , 7'd52 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+261] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+262] = {7'd32 , 8'd72 , 7'd50 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+263] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+264] = {7'd32 , 8'd57 , 7'd47 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+265] = {7'd0  , 8'd7  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+266] = {7'd32 , 8'd44 , 7'd42 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+267] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+268] = {7'd32 , 8'd72 , 7'd39 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+269] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+270] = {7'd32 , 8'd57 , 7'd33 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+271] = {7'd0  , 8'd7  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+272] = {7'd32 , 8'd44 , 7'd29 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+273] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+274] = {7'd32 , 8'd72 , 7'd26 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+275] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+276] = {7'd32 , 8'd57 , 7'd25 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+277] = {7'd0  , 8'd7  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+278] = {7'd32 , 8'd44 , 7'd24 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+279] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+280] = {7'd32 , 8'd72 , 7'd21 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+281] = {7'd0  , 8'd8  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+282] = {7'd32 , 8'd57 , 7'd17 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+283] = {7'd0  , 8'd7  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+284] = {7'd32 , 8'd44 , 7'd15 , 2'd0, 2'd0};   //note: 4E
    assign memory[s1+285] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+286] = {7'd0  , 8'd133, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+287] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song
    assign memory[s1+288] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+289] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+290] = {7'd0  , 8'd0  , 7'd0  , 2'd0, 2'd0};   

    assign memory[s2+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s2+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+79 ] = {7'd0  , 8'd79 , 7'd0  , 2'd0, 2'd0};
    assign memory[s2+80 ] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song
    
    assign memory[s3+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s3+1  ] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+2  ] = {7'd31 , 8'd192, 7'd65 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+3  ] = {7'd31 , 8'd192, 7'd65 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+4  ] = {7'd27 , 8'd192, 7'd65 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+5  ] = {7'd27 , 8'd192, 7'd65 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+6  ] = {7'd27 , 8'd192, 7'd65 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+7  ] = {7'd31 , 8'd192, 7'd65 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+8  ] = {7'd27 , 8'd192, 7'd65 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+9  ] = {7'd31 , 8'd192, 7'd65 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+16 ] = {7'd0  , 8'd6  , 7'd0  , 2'd0, 2'd0};
    assign memory[s3+17 ] = {7'd27 , 8'd188, 7'd79 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+18 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+19 ] = {7'd27 , 8'd188, 7'd79 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+20 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+21 ] = {7'd29 , 8'd188, 7'd79 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s3+22 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+23 ] = {7'd27 , 8'd188, 7'd79 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+24 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+25 ] = {7'd27 , 8'd188, 7'd79 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+26 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+27 ] = {7'd27 , 8'd188, 7'd79 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+28 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+29 ] = {7'd29 , 8'd188, 7'd79 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s3+30 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+31 ] = {7'd27 , 8'd96 , 7'd79 , 2'd0, 2'd0};   //note: 3B
    assign memory[s3+32 ] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+49 ] = {7'd0  , 8'd144, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+50 ] = {7'd28 , 8'd192, 7'd88 , 2'd0, 2'd0};   //note: 4C
    assign memory[s3+51 ] = {7'd29 , 8'd192, 7'd88 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s3+52 ] = {7'd31 , 8'd192, 7'd88 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+53 ] = {7'd28 , 8'd192, 7'd88 , 2'd0, 2'd0};   //note: 4C
    assign memory[s3+54 ] = {7'd29 , 8'd192, 7'd88 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s3+55 ] = {7'd28 , 8'd192, 7'd88 , 2'd0, 2'd0};   //note: 4C
    assign memory[s3+56 ] = {7'd31 , 8'd192, 7'd88 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+57 ] = {7'd28 , 8'd192, 7'd88 , 2'd0, 2'd0};   //note: 4C
    assign memory[s3+58 ] = {7'd33 , 8'd192, 7'd73 , 2'd0, 2'd0};   //note: 4F
    assign memory[s3+59 ] = {7'd33 , 8'd192, 7'd82 , 2'd0, 2'd0};   //note: 4F
    assign memory[s3+60 ] = {7'd35 , 8'd192, 7'd92 , 2'd0, 2'd0};   //note: 4G
    assign memory[s3+61 ] = {7'd36 , 8'd192, 7'd101, 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s3+62 ] = {7'd33 , 8'd192, 7'd98 , 2'd0, 2'd0};   //note: 4F
    assign memory[s3+63 ] = {7'd31 , 8'd192, 7'd95 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s3+64 ] = {7'd29 , 8'd255, 7'd92 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s3+65 ] = {7'd29 , 8'd129, 7'd92 , 2'd0, 2'd0};
    assign memory[s3+66 ] = {7'd29 , 8'd255, 7'd88 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s3+67 ] = {7'd29 , 8'd129, 7'd88 , 2'd0, 2'd0};
    assign memory[s3+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+79 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+80 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+81 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+82 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+83 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+84 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+85 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+86 ] = {7'd0  , 8'd210, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+87 ] = {7'd39 , 8'd96 , 7'd93 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+88 ] = {7'd39 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+89 ] = {7'd39 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+90 ] = {7'd39 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+91 ] = {7'd39 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+92 ] = {7'd39 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+93 ] = {7'd39 , 8'd96 , 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+94 ] = {7'd39 , 8'd255, 7'd88 , 2'd0, 2'd0};   //note: 4B
    assign memory[s3+95 ] = {7'd39 , 8'd225, 7'd88 , 2'd0, 2'd0};
    assign memory[s3+96 ] = {7'd0  , 8'd2  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+97 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+98 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+99 ] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song


endmodule							
