module sine_rom (
    input clk,
	output reg [15:0] dout,
	input [11:0] addr
    );
	
	wire [15:0] memory [4095:0];

	always @(posedge clk) begin
	    dout = memory[addr];
    end
    
    assign memory[   0] = 16'd16384;
    assign memory[   1] = 16'd16409;
    assign memory[   2] = 16'd16434;
    assign memory[   3] = 16'd16459;
    assign memory[   4] = 16'd16484;
    assign memory[   5] = 16'd16509;
    assign memory[   6] = 16'd16534;
    assign memory[   7] = 16'd16559;
    assign memory[   8] = 16'd16585;
    assign memory[   9] = 16'd16610;
    assign memory[  10] = 16'd16635;
    assign memory[  11] = 16'd16660;
    assign memory[  12] = 16'd16685;
    assign memory[  13] = 16'd16710;
    assign memory[  14] = 16'd16735;
    assign memory[  15] = 16'd16760;
    assign memory[  16] = 16'd16786;
    assign memory[  17] = 16'd16811;
    assign memory[  18] = 16'd16836;
    assign memory[  19] = 16'd16861;
    assign memory[  20] = 16'd16886;
    assign memory[  21] = 16'd16911;
    assign memory[  22] = 16'd16936;
    assign memory[  23] = 16'd16961;
    assign memory[  24] = 16'd16987;
    assign memory[  25] = 16'd17012;
    assign memory[  26] = 16'd17037;
    assign memory[  27] = 16'd17062;
    assign memory[  28] = 16'd17087;
    assign memory[  29] = 16'd17112;
    assign memory[  30] = 16'd17137;
    assign memory[  31] = 16'd17162;
    assign memory[  32] = 16'd17187;
    assign memory[  33] = 16'd17213;
    assign memory[  34] = 16'd17238;
    assign memory[  35] = 16'd17263;
    assign memory[  36] = 16'd17288;
    assign memory[  37] = 16'd17313;
    assign memory[  38] = 16'd17338;
    assign memory[  39] = 16'd17363;
    assign memory[  40] = 16'd17388;
    assign memory[  41] = 16'd17413;
    assign memory[  42] = 16'd17438;
    assign memory[  43] = 16'd17463;
    assign memory[  44] = 16'd17489;
    assign memory[  45] = 16'd17514;
    assign memory[  46] = 16'd17539;
    assign memory[  47] = 16'd17564;
    assign memory[  48] = 16'd17589;
    assign memory[  49] = 16'd17614;
    assign memory[  50] = 16'd17639;
    assign memory[  51] = 16'd17664;
    assign memory[  52] = 16'd17689;
    assign memory[  53] = 16'd17714;
    assign memory[  54] = 16'd17739;
    assign memory[  55] = 16'd17764;
    assign memory[  56] = 16'd17789;
    assign memory[  57] = 16'd17814;
    assign memory[  58] = 16'd17839;
    assign memory[  59] = 16'd17864;
    assign memory[  60] = 16'd17889;
    assign memory[  61] = 16'd17914;
    assign memory[  62] = 16'd17939;
    assign memory[  63] = 16'd17964;
    assign memory[  64] = 16'd17989;
    assign memory[  65] = 16'd18014;
    assign memory[  66] = 16'd18039;
    assign memory[  67] = 16'd18064;
    assign memory[  68] = 16'd18089;
    assign memory[  69] = 16'd18114;
    assign memory[  70] = 16'd18139;
    assign memory[  71] = 16'd18164;
    assign memory[  72] = 16'd18189;
    assign memory[  73] = 16'd18214;
    assign memory[  74] = 16'd18239;
    assign memory[  75] = 16'd18264;
    assign memory[  76] = 16'd18289;
    assign memory[  77] = 16'd18314;
    assign memory[  78] = 16'd18339;
    assign memory[  79] = 16'd18364;
    assign memory[  80] = 16'd18389;
    assign memory[  81] = 16'd18414;
    assign memory[  82] = 16'd18439;
    assign memory[  83] = 16'd18464;
    assign memory[  84] = 16'd18489;
    assign memory[  85] = 16'd18514;
    assign memory[  86] = 16'd18539;
    assign memory[  87] = 16'd18564;
    assign memory[  88] = 16'd18588;
    assign memory[  89] = 16'd18613;
    assign memory[  90] = 16'd18638;
    assign memory[  91] = 16'd18663;
    assign memory[  92] = 16'd18688;
    assign memory[  93] = 16'd18713;
    assign memory[  94] = 16'd18738;
    assign memory[  95] = 16'd18763;
    assign memory[  96] = 16'd18788;
    assign memory[  97] = 16'd18812;
    assign memory[  98] = 16'd18837;
    assign memory[  99] = 16'd18862;
    assign memory[ 100] = 16'd18887;
    assign memory[ 101] = 16'd18912;
    assign memory[ 102] = 16'd18937;
    assign memory[ 103] = 16'd18961;
    assign memory[ 104] = 16'd18986;
    assign memory[ 105] = 16'd19011;
    assign memory[ 106] = 16'd19036;
    assign memory[ 107] = 16'd19061;
    assign memory[ 108] = 16'd19085;
    assign memory[ 109] = 16'd19110;
    assign memory[ 110] = 16'd19135;
    assign memory[ 111] = 16'd19160;
    assign memory[ 112] = 16'd19185;
    assign memory[ 113] = 16'd19209;
    assign memory[ 114] = 16'd19234;
    assign memory[ 115] = 16'd19259;
    assign memory[ 116] = 16'd19284;
    assign memory[ 117] = 16'd19308;
    assign memory[ 118] = 16'd19333;
    assign memory[ 119] = 16'd19358;
    assign memory[ 120] = 16'd19382;
    assign memory[ 121] = 16'd19407;
    assign memory[ 122] = 16'd19432;
    assign memory[ 123] = 16'd19457;
    assign memory[ 124] = 16'd19481;
    assign memory[ 125] = 16'd19506;
    assign memory[ 126] = 16'd19531;
    assign memory[ 127] = 16'd19555;
    assign memory[ 128] = 16'd19580;
    assign memory[ 129] = 16'd19605;
    assign memory[ 130] = 16'd19629;
    assign memory[ 131] = 16'd19654;
    assign memory[ 132] = 16'd19678;
    assign memory[ 133] = 16'd19703;
    assign memory[ 134] = 16'd19728;
    assign memory[ 135] = 16'd19752;
    assign memory[ 136] = 16'd19777;
    assign memory[ 137] = 16'd19801;
    assign memory[ 138] = 16'd19826;
    assign memory[ 139] = 16'd19851;
    assign memory[ 140] = 16'd19875;
    assign memory[ 141] = 16'd19900;
    assign memory[ 142] = 16'd19924;
    assign memory[ 143] = 16'd19949;
    assign memory[ 144] = 16'd19973;
    assign memory[ 145] = 16'd19998;
    assign memory[ 146] = 16'd20022;
    assign memory[ 147] = 16'd20047;
    assign memory[ 148] = 16'd20071;
    assign memory[ 149] = 16'd20096;
    assign memory[ 150] = 16'd20120;
    assign memory[ 151] = 16'd20145;
    assign memory[ 152] = 16'd20169;
    assign memory[ 153] = 16'd20194;
    assign memory[ 154] = 16'd20218;
    assign memory[ 155] = 16'd20242;
    assign memory[ 156] = 16'd20267;
    assign memory[ 157] = 16'd20291;
    assign memory[ 158] = 16'd20316;
    assign memory[ 159] = 16'd20340;
    assign memory[ 160] = 16'd20364;
    assign memory[ 161] = 16'd20389;
    assign memory[ 162] = 16'd20413;
    assign memory[ 163] = 16'd20438;
    assign memory[ 164] = 16'd20462;
    assign memory[ 165] = 16'd20486;
    assign memory[ 166] = 16'd20511;
    assign memory[ 167] = 16'd20535;
    assign memory[ 168] = 16'd20559;
    assign memory[ 169] = 16'd20584;
    assign memory[ 170] = 16'd20608;
    assign memory[ 171] = 16'd20632;
    assign memory[ 172] = 16'd20656;
    assign memory[ 173] = 16'd20681;
    assign memory[ 174] = 16'd20705;
    assign memory[ 175] = 16'd20729;
    assign memory[ 176] = 16'd20753;
    assign memory[ 177] = 16'd20778;
    assign memory[ 178] = 16'd20802;
    assign memory[ 179] = 16'd20826;
    assign memory[ 180] = 16'd20850;
    assign memory[ 181] = 16'd20874;
    assign memory[ 182] = 16'd20898;
    assign memory[ 183] = 16'd20923;
    assign memory[ 184] = 16'd20947;
    assign memory[ 185] = 16'd20971;
    assign memory[ 186] = 16'd20995;
    assign memory[ 187] = 16'd21019;
    assign memory[ 188] = 16'd21043;
    assign memory[ 189] = 16'd21067;
    assign memory[ 190] = 16'd21091;
    assign memory[ 191] = 16'd21115;
    assign memory[ 192] = 16'd21140;
    assign memory[ 193] = 16'd21164;
    assign memory[ 194] = 16'd21188;
    assign memory[ 195] = 16'd21212;
    assign memory[ 196] = 16'd21236;
    assign memory[ 197] = 16'd21260;
    assign memory[ 198] = 16'd21284;
    assign memory[ 199] = 16'd21308;
    assign memory[ 200] = 16'd21332;
    assign memory[ 201] = 16'd21356;
    assign memory[ 202] = 16'd21379;
    assign memory[ 203] = 16'd21403;
    assign memory[ 204] = 16'd21427;
    assign memory[ 205] = 16'd21451;
    assign memory[ 206] = 16'd21475;
    assign memory[ 207] = 16'd21499;
    assign memory[ 208] = 16'd21523;
    assign memory[ 209] = 16'd21547;
    assign memory[ 210] = 16'd21571;
    assign memory[ 211] = 16'd21594;
    assign memory[ 212] = 16'd21618;
    assign memory[ 213] = 16'd21642;
    assign memory[ 214] = 16'd21666;
    assign memory[ 215] = 16'd21690;
    assign memory[ 216] = 16'd21713;
    assign memory[ 217] = 16'd21737;
    assign memory[ 218] = 16'd21761;
    assign memory[ 219] = 16'd21785;
    assign memory[ 220] = 16'd21808;
    assign memory[ 221] = 16'd21832;
    assign memory[ 222] = 16'd21856;
    assign memory[ 223] = 16'd21879;
    assign memory[ 224] = 16'd21903;
    assign memory[ 225] = 16'd21927;
    assign memory[ 226] = 16'd21950;
    assign memory[ 227] = 16'd21974;
    assign memory[ 228] = 16'd21998;
    assign memory[ 229] = 16'd22021;
    assign memory[ 230] = 16'd22045;
    assign memory[ 231] = 16'd22068;
    assign memory[ 232] = 16'd22092;
    assign memory[ 233] = 16'd22116;
    assign memory[ 234] = 16'd22139;
    assign memory[ 235] = 16'd22163;
    assign memory[ 236] = 16'd22186;
    assign memory[ 237] = 16'd22210;
    assign memory[ 238] = 16'd22233;
    assign memory[ 239] = 16'd22257;
    assign memory[ 240] = 16'd22280;
    assign memory[ 241] = 16'd22303;
    assign memory[ 242] = 16'd22327;
    assign memory[ 243] = 16'd22350;
    assign memory[ 244] = 16'd22374;
    assign memory[ 245] = 16'd22397;
    assign memory[ 246] = 16'd22420;
    assign memory[ 247] = 16'd22444;
    assign memory[ 248] = 16'd22467;
    assign memory[ 249] = 16'd22490;
    assign memory[ 250] = 16'd22514;
    assign memory[ 251] = 16'd22537;
    assign memory[ 252] = 16'd22560;
    assign memory[ 253] = 16'd22584;
    assign memory[ 254] = 16'd22607;
    assign memory[ 255] = 16'd22630;
    assign memory[ 256] = 16'd22653;
    assign memory[ 257] = 16'd22677;
    assign memory[ 258] = 16'd22700;
    assign memory[ 259] = 16'd22723;
    assign memory[ 260] = 16'd22746;
    assign memory[ 261] = 16'd22769;
    assign memory[ 262] = 16'd22792;
    assign memory[ 263] = 16'd22816;
    assign memory[ 264] = 16'd22839;
    assign memory[ 265] = 16'd22862;
    assign memory[ 266] = 16'd22885;
    assign memory[ 267] = 16'd22908;
    assign memory[ 268] = 16'd22931;
    assign memory[ 269] = 16'd22954;
    assign memory[ 270] = 16'd22977;
    assign memory[ 271] = 16'd23000;
    assign memory[ 272] = 16'd23023;
    assign memory[ 273] = 16'd23046;
    assign memory[ 274] = 16'd23069;
    assign memory[ 275] = 16'd23092;
    assign memory[ 276] = 16'd23115;
    assign memory[ 277] = 16'd23138;
    assign memory[ 278] = 16'd23161;
    assign memory[ 279] = 16'd23183;
    assign memory[ 280] = 16'd23206;
    assign memory[ 281] = 16'd23229;
    assign memory[ 282] = 16'd23252;
    assign memory[ 283] = 16'd23275;
    assign memory[ 284] = 16'd23298;
    assign memory[ 285] = 16'd23320;
    assign memory[ 286] = 16'd23343;
    assign memory[ 287] = 16'd23366;
    assign memory[ 288] = 16'd23389;
    assign memory[ 289] = 16'd23411;
    assign memory[ 290] = 16'd23434;
    assign memory[ 291] = 16'd23457;
    assign memory[ 292] = 16'd23479;
    assign memory[ 293] = 16'd23502;
    assign memory[ 294] = 16'd23525;
    assign memory[ 295] = 16'd23547;
    assign memory[ 296] = 16'd23570;
    assign memory[ 297] = 16'd23592;
    assign memory[ 298] = 16'd23615;
    assign memory[ 299] = 16'd23637;
    assign memory[ 300] = 16'd23660;
    assign memory[ 301] = 16'd23683;
    assign memory[ 302] = 16'd23705;
    assign memory[ 303] = 16'd23727;
    assign memory[ 304] = 16'd23750;
    assign memory[ 305] = 16'd23772;
    assign memory[ 306] = 16'd23795;
    assign memory[ 307] = 16'd23817;
    assign memory[ 308] = 16'd23840;
    assign memory[ 309] = 16'd23862;
    assign memory[ 310] = 16'd23884;
    assign memory[ 311] = 16'd23907;
    assign memory[ 312] = 16'd23929;
    assign memory[ 313] = 16'd23951;
    assign memory[ 314] = 16'd23974;
    assign memory[ 315] = 16'd23996;
    assign memory[ 316] = 16'd24018;
    assign memory[ 317] = 16'd24040;
    assign memory[ 318] = 16'd24062;
    assign memory[ 319] = 16'd24085;
    assign memory[ 320] = 16'd24107;
    assign memory[ 321] = 16'd24129;
    assign memory[ 322] = 16'd24151;
    assign memory[ 323] = 16'd24173;
    assign memory[ 324] = 16'd24195;
    assign memory[ 325] = 16'd24217;
    assign memory[ 326] = 16'd24240;
    assign memory[ 327] = 16'd24262;
    assign memory[ 328] = 16'd24284;
    assign memory[ 329] = 16'd24306;
    assign memory[ 330] = 16'd24328;
    assign memory[ 331] = 16'd24350;
    assign memory[ 332] = 16'd24372;
    assign memory[ 333] = 16'd24393;
    assign memory[ 334] = 16'd24415;
    assign memory[ 335] = 16'd24437;
    assign memory[ 336] = 16'd24459;
    assign memory[ 337] = 16'd24481;
    assign memory[ 338] = 16'd24503;
    assign memory[ 339] = 16'd24525;
    assign memory[ 340] = 16'd24546;
    assign memory[ 341] = 16'd24568;
    assign memory[ 342] = 16'd24590;
    assign memory[ 343] = 16'd24612;
    assign memory[ 344] = 16'd24633;
    assign memory[ 345] = 16'd24655;
    assign memory[ 346] = 16'd24677;
    assign memory[ 347] = 16'd24699;
    assign memory[ 348] = 16'd24720;
    assign memory[ 349] = 16'd24742;
    assign memory[ 350] = 16'd24763;
    assign memory[ 351] = 16'd24785;
    assign memory[ 352] = 16'd24807;
    assign memory[ 353] = 16'd24828;
    assign memory[ 354] = 16'd24850;
    assign memory[ 355] = 16'd24871;
    assign memory[ 356] = 16'd24893;
    assign memory[ 357] = 16'd24914;
    assign memory[ 358] = 16'd24936;
    assign memory[ 359] = 16'd24957;
    assign memory[ 360] = 16'd24978;
    assign memory[ 361] = 16'd25000;
    assign memory[ 362] = 16'd25021;
    assign memory[ 363] = 16'd25042;
    assign memory[ 364] = 16'd25064;
    assign memory[ 365] = 16'd25085;
    assign memory[ 366] = 16'd25106;
    assign memory[ 367] = 16'd25128;
    assign memory[ 368] = 16'd25149;
    assign memory[ 369] = 16'd25170;
    assign memory[ 370] = 16'd25191;
    assign memory[ 371] = 16'd25213;
    assign memory[ 372] = 16'd25234;
    assign memory[ 373] = 16'd25255;
    assign memory[ 374] = 16'd25276;
    assign memory[ 375] = 16'd25297;
    assign memory[ 376] = 16'd25318;
    assign memory[ 377] = 16'd25339;
    assign memory[ 378] = 16'd25360;
    assign memory[ 379] = 16'd25381;
    assign memory[ 380] = 16'd25402;
    assign memory[ 381] = 16'd25423;
    assign memory[ 382] = 16'd25444;
    assign memory[ 383] = 16'd25465;
    assign memory[ 384] = 16'd25486;
    assign memory[ 385] = 16'd25507;
    assign memory[ 386] = 16'd25528;
    assign memory[ 387] = 16'd25549;
    assign memory[ 388] = 16'd25569;
    assign memory[ 389] = 16'd25590;
    assign memory[ 390] = 16'd25611;
    assign memory[ 391] = 16'd25632;
    assign memory[ 392] = 16'd25652;
    assign memory[ 393] = 16'd25673;
    assign memory[ 394] = 16'd25694;
    assign memory[ 395] = 16'd25715;
    assign memory[ 396] = 16'd25735;
    assign memory[ 397] = 16'd25756;
    assign memory[ 398] = 16'd25776;
    assign memory[ 399] = 16'd25797;
    assign memory[ 400] = 16'd25818;
    assign memory[ 401] = 16'd25838;
    assign memory[ 402] = 16'd25859;
    assign memory[ 403] = 16'd25879;
    assign memory[ 404] = 16'd25900;
    assign memory[ 405] = 16'd25920;
    assign memory[ 406] = 16'd25940;
    assign memory[ 407] = 16'd25961;
    assign memory[ 408] = 16'd25981;
    assign memory[ 409] = 16'd26002;
    assign memory[ 410] = 16'd26022;
    assign memory[ 411] = 16'd26042;
    assign memory[ 412] = 16'd26063;
    assign memory[ 413] = 16'd26083;
    assign memory[ 414] = 16'd26103;
    assign memory[ 415] = 16'd26123;
    assign memory[ 416] = 16'd26143;
    assign memory[ 417] = 16'd26164;
    assign memory[ 418] = 16'd26184;
    assign memory[ 419] = 16'd26204;
    assign memory[ 420] = 16'd26224;
    assign memory[ 421] = 16'd26244;
    assign memory[ 422] = 16'd26264;
    assign memory[ 423] = 16'd26284;
    assign memory[ 424] = 16'd26304;
    assign memory[ 425] = 16'd26324;
    assign memory[ 426] = 16'd26344;
    assign memory[ 427] = 16'd26364;
    assign memory[ 428] = 16'd26384;
    assign memory[ 429] = 16'd26404;
    assign memory[ 430] = 16'd26424;
    assign memory[ 431] = 16'd26444;
    assign memory[ 432] = 16'd26463;
    assign memory[ 433] = 16'd26483;
    assign memory[ 434] = 16'd26503;
    assign memory[ 435] = 16'd26523;
    assign memory[ 436] = 16'd26543;
    assign memory[ 437] = 16'd26562;
    assign memory[ 438] = 16'd26582;
    assign memory[ 439] = 16'd26602;
    assign memory[ 440] = 16'd26621;
    assign memory[ 441] = 16'd26641;
    assign memory[ 442] = 16'd26660;
    assign memory[ 443] = 16'd26680;
    assign memory[ 444] = 16'd26699;
    assign memory[ 445] = 16'd26719;
    assign memory[ 446] = 16'd26738;
    assign memory[ 447] = 16'd26758;
    assign memory[ 448] = 16'd26777;
    assign memory[ 449] = 16'd26797;
    assign memory[ 450] = 16'd26816;
    assign memory[ 451] = 16'd26836;
    assign memory[ 452] = 16'd26855;
    assign memory[ 453] = 16'd26874;
    assign memory[ 454] = 16'd26894;
    assign memory[ 455] = 16'd26913;
    assign memory[ 456] = 16'd26932;
    assign memory[ 457] = 16'd26951;
    assign memory[ 458] = 16'd26970;
    assign memory[ 459] = 16'd26990;
    assign memory[ 460] = 16'd27009;
    assign memory[ 461] = 16'd27028;
    assign memory[ 462] = 16'd27047;
    assign memory[ 463] = 16'd27066;
    assign memory[ 464] = 16'd27085;
    assign memory[ 465] = 16'd27104;
    assign memory[ 466] = 16'd27123;
    assign memory[ 467] = 16'd27142;
    assign memory[ 468] = 16'd27161;
    assign memory[ 469] = 16'd27180;
    assign memory[ 470] = 16'd27199;
    assign memory[ 471] = 16'd27218;
    assign memory[ 472] = 16'd27237;
    assign memory[ 473] = 16'd27255;
    assign memory[ 474] = 16'd27274;
    assign memory[ 475] = 16'd27293;
    assign memory[ 476] = 16'd27312;
    assign memory[ 477] = 16'd27330;
    assign memory[ 478] = 16'd27349;
    assign memory[ 479] = 16'd27368;
    assign memory[ 480] = 16'd27386;
    assign memory[ 481] = 16'd27405;
    assign memory[ 482] = 16'd27424;
    assign memory[ 483] = 16'd27442;
    assign memory[ 484] = 16'd27461;
    assign memory[ 485] = 16'd27479;
    assign memory[ 486] = 16'd27498;
    assign memory[ 487] = 16'd27516;
    assign memory[ 488] = 16'd27534;
    assign memory[ 489] = 16'd27553;
    assign memory[ 490] = 16'd27571;
    assign memory[ 491] = 16'd27590;
    assign memory[ 492] = 16'd27608;
    assign memory[ 493] = 16'd27626;
    assign memory[ 494] = 16'd27644;
    assign memory[ 495] = 16'd27663;
    assign memory[ 496] = 16'd27681;
    assign memory[ 497] = 16'd27699;
    assign memory[ 498] = 16'd27717;
    assign memory[ 499] = 16'd27735;
    assign memory[ 500] = 16'd27754;
    assign memory[ 501] = 16'd27772;
    assign memory[ 502] = 16'd27790;
    assign memory[ 503] = 16'd27808;
    assign memory[ 504] = 16'd27826;
    assign memory[ 505] = 16'd27844;
    assign memory[ 506] = 16'd27862;
    assign memory[ 507] = 16'd27880;
    assign memory[ 508] = 16'd27897;
    assign memory[ 509] = 16'd27915;
    assign memory[ 510] = 16'd27933;
    assign memory[ 511] = 16'd27951;
    assign memory[ 512] = 16'd27969;
    assign memory[ 513] = 16'd27986;
    assign memory[ 514] = 16'd28004;
    assign memory[ 515] = 16'd28022;
    assign memory[ 516] = 16'd28040;
    assign memory[ 517] = 16'd28057;
    assign memory[ 518] = 16'd28075;
    assign memory[ 519] = 16'd28092;
    assign memory[ 520] = 16'd28110;
    assign memory[ 521] = 16'd28128;
    assign memory[ 522] = 16'd28145;
    assign memory[ 523] = 16'd28163;
    assign memory[ 524] = 16'd28180;
    assign memory[ 525] = 16'd28197;
    assign memory[ 526] = 16'd28215;
    assign memory[ 527] = 16'd28232;
    assign memory[ 528] = 16'd28250;
    assign memory[ 529] = 16'd28267;
    assign memory[ 530] = 16'd28284;
    assign memory[ 531] = 16'd28301;
    assign memory[ 532] = 16'd28319;
    assign memory[ 533] = 16'd28336;
    assign memory[ 534] = 16'd28353;
    assign memory[ 535] = 16'd28370;
    assign memory[ 536] = 16'd28387;
    assign memory[ 537] = 16'd28404;
    assign memory[ 538] = 16'd28421;
    assign memory[ 539] = 16'd28438;
    assign memory[ 540] = 16'd28456;
    assign memory[ 541] = 16'd28472;
    assign memory[ 542] = 16'd28489;
    assign memory[ 543] = 16'd28506;
    assign memory[ 544] = 16'd28523;
    assign memory[ 545] = 16'd28540;
    assign memory[ 546] = 16'd28557;
    assign memory[ 547] = 16'd28574;
    assign memory[ 548] = 16'd28591;
    assign memory[ 549] = 16'd28607;
    assign memory[ 550] = 16'd28624;
    assign memory[ 551] = 16'd28641;
    assign memory[ 552] = 16'd28657;
    assign memory[ 553] = 16'd28674;
    assign memory[ 554] = 16'd28691;
    assign memory[ 555] = 16'd28707;
    assign memory[ 556] = 16'd28724;
    assign memory[ 557] = 16'd28740;
    assign memory[ 558] = 16'd28757;
    assign memory[ 559] = 16'd28773;
    assign memory[ 560] = 16'd28790;
    assign memory[ 561] = 16'd28806;
    assign memory[ 562] = 16'd28822;
    assign memory[ 563] = 16'd28839;
    assign memory[ 564] = 16'd28855;
    assign memory[ 565] = 16'd28871;
    assign memory[ 566] = 16'd28888;
    assign memory[ 567] = 16'd28904;
    assign memory[ 568] = 16'd28920;
    assign memory[ 569] = 16'd28936;
    assign memory[ 570] = 16'd28952;
    assign memory[ 571] = 16'd28968;
    assign memory[ 572] = 16'd28984;
    assign memory[ 573] = 16'd29001;
    assign memory[ 574] = 16'd29017;
    assign memory[ 575] = 16'd29033;
    assign memory[ 576] = 16'd29049;
    assign memory[ 577] = 16'd29064;
    assign memory[ 578] = 16'd29080;
    assign memory[ 579] = 16'd29096;
    assign memory[ 580] = 16'd29112;
    assign memory[ 581] = 16'd29128;
    assign memory[ 582] = 16'd29144;
    assign memory[ 583] = 16'd29159;
    assign memory[ 584] = 16'd29175;
    assign memory[ 585] = 16'd29191;
    assign memory[ 586] = 16'd29206;
    assign memory[ 587] = 16'd29222;
    assign memory[ 588] = 16'd29238;
    assign memory[ 589] = 16'd29253;
    assign memory[ 590] = 16'd29269;
    assign memory[ 591] = 16'd29284;
    assign memory[ 592] = 16'd29300;
    assign memory[ 593] = 16'd29315;
    assign memory[ 594] = 16'd29331;
    assign memory[ 595] = 16'd29346;
    assign memory[ 596] = 16'd29361;
    assign memory[ 597] = 16'd29377;
    assign memory[ 598] = 16'd29392;
    assign memory[ 599] = 16'd29407;
    assign memory[ 600] = 16'd29422;
    assign memory[ 601] = 16'd29438;
    assign memory[ 602] = 16'd29453;
    assign memory[ 603] = 16'd29468;
    assign memory[ 604] = 16'd29483;
    assign memory[ 605] = 16'd29498;
    assign memory[ 606] = 16'd29513;
    assign memory[ 607] = 16'd29528;
    assign memory[ 608] = 16'd29543;
    assign memory[ 609] = 16'd29558;
    assign memory[ 610] = 16'd29573;
    assign memory[ 611] = 16'd29588;
    assign memory[ 612] = 16'd29603;
    assign memory[ 613] = 16'd29618;
    assign memory[ 614] = 16'd29633;
    assign memory[ 615] = 16'd29647;
    assign memory[ 616] = 16'd29662;
    assign memory[ 617] = 16'd29677;
    assign memory[ 618] = 16'd29691;
    assign memory[ 619] = 16'd29706;
    assign memory[ 620] = 16'd29721;
    assign memory[ 621] = 16'd29735;
    assign memory[ 622] = 16'd29750;
    assign memory[ 623] = 16'd29764;
    assign memory[ 624] = 16'd29779;
    assign memory[ 625] = 16'd29793;
    assign memory[ 626] = 16'd29808;
    assign memory[ 627] = 16'd29822;
    assign memory[ 628] = 16'd29836;
    assign memory[ 629] = 16'd29851;
    assign memory[ 630] = 16'd29865;
    assign memory[ 631] = 16'd29879;
    assign memory[ 632] = 16'd29894;
    assign memory[ 633] = 16'd29908;
    assign memory[ 634] = 16'd29922;
    assign memory[ 635] = 16'd29936;
    assign memory[ 636] = 16'd29950;
    assign memory[ 637] = 16'd29964;
    assign memory[ 638] = 16'd29978;
    assign memory[ 639] = 16'd29992;
    assign memory[ 640] = 16'd30006;
    assign memory[ 641] = 16'd30020;
    assign memory[ 642] = 16'd30034;
    assign memory[ 643] = 16'd30048;
    assign memory[ 644] = 16'd30062;
    assign memory[ 645] = 16'd30076;
    assign memory[ 646] = 16'd30089;
    assign memory[ 647] = 16'd30103;
    assign memory[ 648] = 16'd30117;
    assign memory[ 649] = 16'd30131;
    assign memory[ 650] = 16'd30144;
    assign memory[ 651] = 16'd30158;
    assign memory[ 652] = 16'd30172;
    assign memory[ 653] = 16'd30185;
    assign memory[ 654] = 16'd30199;
    assign memory[ 655] = 16'd30212;
    assign memory[ 656] = 16'd30226;
    assign memory[ 657] = 16'd30239;
    assign memory[ 658] = 16'd30252;
    assign memory[ 659] = 16'd30266;
    assign memory[ 660] = 16'd30279;
    assign memory[ 661] = 16'd30292;
    assign memory[ 662] = 16'd30306;
    assign memory[ 663] = 16'd30319;
    assign memory[ 664] = 16'd30332;
    assign memory[ 665] = 16'd30345;
    assign memory[ 666] = 16'd30358;
    assign memory[ 667] = 16'd30372;
    assign memory[ 668] = 16'd30385;
    assign memory[ 669] = 16'd30398;
    assign memory[ 670] = 16'd30411;
    assign memory[ 671] = 16'd30424;
    assign memory[ 672] = 16'd30437;
    assign memory[ 673] = 16'd30449;
    assign memory[ 674] = 16'd30462;
    assign memory[ 675] = 16'd30475;
    assign memory[ 676] = 16'd30488;
    assign memory[ 677] = 16'd30501;
    assign memory[ 678] = 16'd30513;
    assign memory[ 679] = 16'd30526;
    assign memory[ 680] = 16'd30539;
    assign memory[ 681] = 16'd30551;
    assign memory[ 682] = 16'd30564;
    assign memory[ 683] = 16'd30577;
    assign memory[ 684] = 16'd30589;
    assign memory[ 685] = 16'd30602;
    assign memory[ 686] = 16'd30614;
    assign memory[ 687] = 16'd30627;
    assign memory[ 688] = 16'd30639;
    assign memory[ 689] = 16'd30651;
    assign memory[ 690] = 16'd30664;
    assign memory[ 691] = 16'd30676;
    assign memory[ 692] = 16'd30688;
    assign memory[ 693] = 16'd30701;
    assign memory[ 694] = 16'd30713;
    assign memory[ 695] = 16'd30725;
    assign memory[ 696] = 16'd30737;
    assign memory[ 697] = 16'd30749;
    assign memory[ 698] = 16'd30761;
    assign memory[ 699] = 16'd30773;
    assign memory[ 700] = 16'd30785;
    assign memory[ 701] = 16'd30797;
    assign memory[ 702] = 16'd30809;
    assign memory[ 703] = 16'd30821;
    assign memory[ 704] = 16'd30833;
    assign memory[ 705] = 16'd30845;
    assign memory[ 706] = 16'd30857;
    assign memory[ 707] = 16'd30868;
    assign memory[ 708] = 16'd30880;
    assign memory[ 709] = 16'd30892;
    assign memory[ 710] = 16'd30903;
    assign memory[ 711] = 16'd30915;
    assign memory[ 712] = 16'd30927;
    assign memory[ 713] = 16'd30938;
    assign memory[ 714] = 16'd30950;
    assign memory[ 715] = 16'd30961;
    assign memory[ 716] = 16'd30973;
    assign memory[ 717] = 16'd30984;
    assign memory[ 718] = 16'd30995;
    assign memory[ 719] = 16'd31007;
    assign memory[ 720] = 16'd31018;
    assign memory[ 721] = 16'd31029;
    assign memory[ 722] = 16'd31041;
    assign memory[ 723] = 16'd31052;
    assign memory[ 724] = 16'd31063;
    assign memory[ 725] = 16'd31074;
    assign memory[ 726] = 16'd31085;
    assign memory[ 727] = 16'd31096;
    assign memory[ 728] = 16'd31107;
    assign memory[ 729] = 16'd31118;
    assign memory[ 730] = 16'd31129;
    assign memory[ 731] = 16'd31140;
    assign memory[ 732] = 16'd31151;
    assign memory[ 733] = 16'd31162;
    assign memory[ 734] = 16'd31173;
    assign memory[ 735] = 16'd31184;
    assign memory[ 736] = 16'd31194;
    assign memory[ 737] = 16'd31205;
    assign memory[ 738] = 16'd31216;
    assign memory[ 739] = 16'd31227;
    assign memory[ 740] = 16'd31237;
    assign memory[ 741] = 16'd31248;
    assign memory[ 742] = 16'd31258;
    assign memory[ 743] = 16'd31269;
    assign memory[ 744] = 16'd31279;
    assign memory[ 745] = 16'd31290;
    assign memory[ 746] = 16'd31300;
    assign memory[ 747] = 16'd31311;
    assign memory[ 748] = 16'd31321;
    assign memory[ 749] = 16'd31331;
    assign memory[ 750] = 16'd31341;
    assign memory[ 751] = 16'd31352;
    assign memory[ 752] = 16'd31362;
    assign memory[ 753] = 16'd31372;
    assign memory[ 754] = 16'd31382;
    assign memory[ 755] = 16'd31392;
    assign memory[ 756] = 16'd31402;
    assign memory[ 757] = 16'd31412;
    assign memory[ 758] = 16'd31422;
    assign memory[ 759] = 16'd31432;
    assign memory[ 760] = 16'd31442;
    assign memory[ 761] = 16'd31452;
    assign memory[ 762] = 16'd31462;
    assign memory[ 763] = 16'd31472;
    assign memory[ 764] = 16'd31482;
    assign memory[ 765] = 16'd31491;
    assign memory[ 766] = 16'd31501;
    assign memory[ 767] = 16'd31511;
    assign memory[ 768] = 16'd31520;
    assign memory[ 769] = 16'd31530;
    assign memory[ 770] = 16'd31540;
    assign memory[ 771] = 16'd31549;
    assign memory[ 772] = 16'd31559;
    assign memory[ 773] = 16'd31568;
    assign memory[ 774] = 16'd31577;
    assign memory[ 775] = 16'd31587;
    assign memory[ 776] = 16'd31596;
    assign memory[ 777] = 16'd31605;
    assign memory[ 778] = 16'd31615;
    assign memory[ 779] = 16'd31624;
    assign memory[ 780] = 16'd31633;
    assign memory[ 781] = 16'd31642;
    assign memory[ 782] = 16'd31651;
    assign memory[ 783] = 16'd31661;
    assign memory[ 784] = 16'd31670;
    assign memory[ 785] = 16'd31679;
    assign memory[ 786] = 16'd31688;
    assign memory[ 787] = 16'd31697;
    assign memory[ 788] = 16'd31706;
    assign memory[ 789] = 16'd31714;
    assign memory[ 790] = 16'd31723;
    assign memory[ 791] = 16'd31732;
    assign memory[ 792] = 16'd31741;
    assign memory[ 793] = 16'd31750;
    assign memory[ 794] = 16'd31758;
    assign memory[ 795] = 16'd31767;
    assign memory[ 796] = 16'd31776;
    assign memory[ 797] = 16'd31784;
    assign memory[ 798] = 16'd31793;
    assign memory[ 799] = 16'd31801;
    assign memory[ 800] = 16'd31810;
    assign memory[ 801] = 16'd31818;
    assign memory[ 802] = 16'd31827;
    assign memory[ 803] = 16'd31835;
    assign memory[ 804] = 16'd31843;
    assign memory[ 805] = 16'd31852;
    assign memory[ 806] = 16'd31860;
    assign memory[ 807] = 16'd31868;
    assign memory[ 808] = 16'd31876;
    assign memory[ 809] = 16'd31884;
    assign memory[ 810] = 16'd31893;
    assign memory[ 811] = 16'd31901;
    assign memory[ 812] = 16'd31909;
    assign memory[ 813] = 16'd31917;
    assign memory[ 814] = 16'd31925;
    assign memory[ 815] = 16'd31933;
    assign memory[ 816] = 16'd31941;
    assign memory[ 817] = 16'd31948;
    assign memory[ 818] = 16'd31956;
    assign memory[ 819] = 16'd31964;
    assign memory[ 820] = 16'd31972;
    assign memory[ 821] = 16'd31980;
    assign memory[ 822] = 16'd31987;
    assign memory[ 823] = 16'd31995;
    assign memory[ 824] = 16'd32002;
    assign memory[ 825] = 16'd32010;
    assign memory[ 826] = 16'd32018;
    assign memory[ 827] = 16'd32025;
    assign memory[ 828] = 16'd32033;
    assign memory[ 829] = 16'd32040;
    assign memory[ 830] = 16'd32047;
    assign memory[ 831] = 16'd32055;
    assign memory[ 832] = 16'd32062;
    assign memory[ 833] = 16'd32069;
    assign memory[ 834] = 16'd32077;
    assign memory[ 835] = 16'd32084;
    assign memory[ 836] = 16'd32091;
    assign memory[ 837] = 16'd32098;
    assign memory[ 838] = 16'd32105;
    assign memory[ 839] = 16'd32112;
    assign memory[ 840] = 16'd32119;
    assign memory[ 841] = 16'd32126;
    assign memory[ 842] = 16'd32133;
    assign memory[ 843] = 16'd32140;
    assign memory[ 844] = 16'd32147;
    assign memory[ 845] = 16'd32154;
    assign memory[ 846] = 16'd32161;
    assign memory[ 847] = 16'd32167;
    assign memory[ 848] = 16'd32174;
    assign memory[ 849] = 16'd32181;
    assign memory[ 850] = 16'd32187;
    assign memory[ 851] = 16'd32194;
    assign memory[ 852] = 16'd32201;
    assign memory[ 853] = 16'd32207;
    assign memory[ 854] = 16'd32214;
    assign memory[ 855] = 16'd32220;
    assign memory[ 856] = 16'd32226;
    assign memory[ 857] = 16'd32233;
    assign memory[ 858] = 16'd32239;
    assign memory[ 859] = 16'd32245;
    assign memory[ 860] = 16'd32252;
    assign memory[ 861] = 16'd32258;
    assign memory[ 862] = 16'd32264;
    assign memory[ 863] = 16'd32270;
    assign memory[ 864] = 16'd32276;
    assign memory[ 865] = 16'd32283;
    assign memory[ 866] = 16'd32289;
    assign memory[ 867] = 16'd32295;
    assign memory[ 868] = 16'd32301;
    assign memory[ 869] = 16'd32307;
    assign memory[ 870] = 16'd32312;
    assign memory[ 871] = 16'd32318;
    assign memory[ 872] = 16'd32324;
    assign memory[ 873] = 16'd32330;
    assign memory[ 874] = 16'd32336;
    assign memory[ 875] = 16'd32341;
    assign memory[ 876] = 16'd32347;
    assign memory[ 877] = 16'd32353;
    assign memory[ 878] = 16'd32358;
    assign memory[ 879] = 16'd32364;
    assign memory[ 880] = 16'd32369;
    assign memory[ 881] = 16'd32375;
    assign memory[ 882] = 16'd32380;
    assign memory[ 883] = 16'd32386;
    assign memory[ 884] = 16'd32391;
    assign memory[ 885] = 16'd32396;
    assign memory[ 886] = 16'd32402;
    assign memory[ 887] = 16'd32407;
    assign memory[ 888] = 16'd32412;
    assign memory[ 889] = 16'd32417;
    assign memory[ 890] = 16'd32423;
    assign memory[ 891] = 16'd32428;
    assign memory[ 892] = 16'd32433;
    assign memory[ 893] = 16'd32438;
    assign memory[ 894] = 16'd32443;
    assign memory[ 895] = 16'd32448;
    assign memory[ 896] = 16'd32453;
    assign memory[ 897] = 16'd32458;
    assign memory[ 898] = 16'd32462;
    assign memory[ 899] = 16'd32467;
    assign memory[ 900] = 16'd32472;
    assign memory[ 901] = 16'd32477;
    assign memory[ 902] = 16'd32481;
    assign memory[ 903] = 16'd32486;
    assign memory[ 904] = 16'd32491;
    assign memory[ 905] = 16'd32495;
    assign memory[ 906] = 16'd32500;
    assign memory[ 907] = 16'd32504;
    assign memory[ 908] = 16'd32509;
    assign memory[ 909] = 16'd32513;
    assign memory[ 910] = 16'd32518;
    assign memory[ 911] = 16'd32522;
    assign memory[ 912] = 16'd32526;
    assign memory[ 913] = 16'd32531;
    assign memory[ 914] = 16'd32535;
    assign memory[ 915] = 16'd32539;
    assign memory[ 916] = 16'd32543;
    assign memory[ 917] = 16'd32547;
    assign memory[ 918] = 16'd32551;
    assign memory[ 919] = 16'd32555;
    assign memory[ 920] = 16'd32559;
    assign memory[ 921] = 16'd32563;
    assign memory[ 922] = 16'd32567;
    assign memory[ 923] = 16'd32571;
    assign memory[ 924] = 16'd32575;
    assign memory[ 925] = 16'd32579;
    assign memory[ 926] = 16'd32583;
    assign memory[ 927] = 16'd32586;
    assign memory[ 928] = 16'd32590;
    assign memory[ 929] = 16'd32594;
    assign memory[ 930] = 16'd32597;
    assign memory[ 931] = 16'd32601;
    assign memory[ 932] = 16'd32605;
    assign memory[ 933] = 16'd32608;
    assign memory[ 934] = 16'd32612;
    assign memory[ 935] = 16'd32615;
    assign memory[ 936] = 16'd32618;
    assign memory[ 937] = 16'd32622;
    assign memory[ 938] = 16'd32625;
    assign memory[ 939] = 16'd32628;
    assign memory[ 940] = 16'd32632;
    assign memory[ 941] = 16'd32635;
    assign memory[ 942] = 16'd32638;
    assign memory[ 943] = 16'd32641;
    assign memory[ 944] = 16'd32644;
    assign memory[ 945] = 16'd32647;
    assign memory[ 946] = 16'd32650;
    assign memory[ 947] = 16'd32653;
    assign memory[ 948] = 16'd32656;
    assign memory[ 949] = 16'd32659;
    assign memory[ 950] = 16'd32662;
    assign memory[ 951] = 16'd32665;
    assign memory[ 952] = 16'd32668;
    assign memory[ 953] = 16'd32670;
    assign memory[ 954] = 16'd32673;
    assign memory[ 955] = 16'd32676;
    assign memory[ 956] = 16'd32678;
    assign memory[ 957] = 16'd32681;
    assign memory[ 958] = 16'd32684;
    assign memory[ 959] = 16'd32686;
    assign memory[ 960] = 16'd32689;
    assign memory[ 961] = 16'd32691;
    assign memory[ 962] = 16'd32693;
    assign memory[ 963] = 16'd32696;
    assign memory[ 964] = 16'd32698;
    assign memory[ 965] = 16'd32700;
    assign memory[ 966] = 16'd32703;
    assign memory[ 967] = 16'd32705;
    assign memory[ 968] = 16'd32707;
    assign memory[ 969] = 16'd32709;
    assign memory[ 970] = 16'd32711;
    assign memory[ 971] = 16'd32713;
    assign memory[ 972] = 16'd32715;
    assign memory[ 973] = 16'd32717;
    assign memory[ 974] = 16'd32719;
    assign memory[ 975] = 16'd32721;
    assign memory[ 976] = 16'd32723;
    assign memory[ 977] = 16'd32725;
    assign memory[ 978] = 16'd32727;
    assign memory[ 979] = 16'd32728;
    assign memory[ 980] = 16'd32730;
    assign memory[ 981] = 16'd32732;
    assign memory[ 982] = 16'd32734;
    assign memory[ 983] = 16'd32735;
    assign memory[ 984] = 16'd32737;
    assign memory[ 985] = 16'd32738;
    assign memory[ 986] = 16'd32740;
    assign memory[ 987] = 16'd32741;
    assign memory[ 988] = 16'd32743;
    assign memory[ 989] = 16'd32744;
    assign memory[ 990] = 16'd32745;
    assign memory[ 991] = 16'd32747;
    assign memory[ 992] = 16'd32748;
    assign memory[ 993] = 16'd32749;
    assign memory[ 994] = 16'd32750;
    assign memory[ 995] = 16'd32751;
    assign memory[ 996] = 16'd32752;
    assign memory[ 997] = 16'd32753;
    assign memory[ 998] = 16'd32754;
    assign memory[ 999] = 16'd32755;
    assign memory[1000] = 16'd32756;
    assign memory[1001] = 16'd32757;
    assign memory[1002] = 16'd32758;
    assign memory[1003] = 16'd32759;
    assign memory[1004] = 16'd32760;
    assign memory[1005] = 16'd32761;
    assign memory[1006] = 16'd32761;
    assign memory[1007] = 16'd32762;
    assign memory[1008] = 16'd32763;
    assign memory[1009] = 16'd32763;
    assign memory[1010] = 16'd32764;
    assign memory[1011] = 16'd32764;
    assign memory[1012] = 16'd32765;
    assign memory[1013] = 16'd32765;
    assign memory[1014] = 16'd32766;
    assign memory[1015] = 16'd32766;
    assign memory[1016] = 16'd32766;
    assign memory[1017] = 16'd32767;
    assign memory[1018] = 16'd32767;
    assign memory[1019] = 16'd32767;
    assign memory[1020] = 16'd32767;
    assign memory[1021] = 16'd32767;
    assign memory[1022] = 16'd32767;
    assign memory[1023] = 16'd32767;
    assign memory[1024] = 16'd32767;
    assign memory[1025] = 16'd32767;
    assign memory[1026] = 16'd32767;
    assign memory[1027] = 16'd32767;
    assign memory[1028] = 16'd32767;
    assign memory[1029] = 16'd32767;
    assign memory[1030] = 16'd32767;
    assign memory[1031] = 16'd32767;
    assign memory[1032] = 16'd32766;
    assign memory[1033] = 16'd32766;
    assign memory[1034] = 16'd32766;
    assign memory[1035] = 16'd32765;
    assign memory[1036] = 16'd32765;
    assign memory[1037] = 16'd32764;
    assign memory[1038] = 16'd32764;
    assign memory[1039] = 16'd32763;
    assign memory[1040] = 16'd32763;
    assign memory[1041] = 16'd32762;
    assign memory[1042] = 16'd32761;
    assign memory[1043] = 16'd32761;
    assign memory[1044] = 16'd32760;
    assign memory[1045] = 16'd32759;
    assign memory[1046] = 16'd32758;
    assign memory[1047] = 16'd32757;
    assign memory[1048] = 16'd32756;
    assign memory[1049] = 16'd32755;
    assign memory[1050] = 16'd32754;
    assign memory[1051] = 16'd32753;
    assign memory[1052] = 16'd32752;
    assign memory[1053] = 16'd32751;
    assign memory[1054] = 16'd32750;
    assign memory[1055] = 16'd32749;
    assign memory[1056] = 16'd32748;
    assign memory[1057] = 16'd32747;
    assign memory[1058] = 16'd32745;
    assign memory[1059] = 16'd32744;
    assign memory[1060] = 16'd32743;
    assign memory[1061] = 16'd32741;
    assign memory[1062] = 16'd32740;
    assign memory[1063] = 16'd32738;
    assign memory[1064] = 16'd32737;
    assign memory[1065] = 16'd32735;
    assign memory[1066] = 16'd32734;
    assign memory[1067] = 16'd32732;
    assign memory[1068] = 16'd32730;
    assign memory[1069] = 16'd32728;
    assign memory[1070] = 16'd32727;
    assign memory[1071] = 16'd32725;
    assign memory[1072] = 16'd32723;
    assign memory[1073] = 16'd32721;
    assign memory[1074] = 16'd32719;
    assign memory[1075] = 16'd32717;
    assign memory[1076] = 16'd32715;
    assign memory[1077] = 16'd32713;
    assign memory[1078] = 16'd32711;
    assign memory[1079] = 16'd32709;
    assign memory[1080] = 16'd32707;
    assign memory[1081] = 16'd32705;
    assign memory[1082] = 16'd32703;
    assign memory[1083] = 16'd32700;
    assign memory[1084] = 16'd32698;
    assign memory[1085] = 16'd32696;
    assign memory[1086] = 16'd32693;
    assign memory[1087] = 16'd32691;
    assign memory[1088] = 16'd32689;
    assign memory[1089] = 16'd32686;
    assign memory[1090] = 16'd32684;
    assign memory[1091] = 16'd32681;
    assign memory[1092] = 16'd32678;
    assign memory[1093] = 16'd32676;
    assign memory[1094] = 16'd32673;
    assign memory[1095] = 16'd32670;
    assign memory[1096] = 16'd32668;
    assign memory[1097] = 16'd32665;
    assign memory[1098] = 16'd32662;
    assign memory[1099] = 16'd32659;
    assign memory[1100] = 16'd32656;
    assign memory[1101] = 16'd32653;
    assign memory[1102] = 16'd32650;
    assign memory[1103] = 16'd32647;
    assign memory[1104] = 16'd32644;
    assign memory[1105] = 16'd32641;
    assign memory[1106] = 16'd32638;
    assign memory[1107] = 16'd32635;
    assign memory[1108] = 16'd32632;
    assign memory[1109] = 16'd32628;
    assign memory[1110] = 16'd32625;
    assign memory[1111] = 16'd32622;
    assign memory[1112] = 16'd32618;
    assign memory[1113] = 16'd32615;
    assign memory[1114] = 16'd32612;
    assign memory[1115] = 16'd32608;
    assign memory[1116] = 16'd32605;
    assign memory[1117] = 16'd32601;
    assign memory[1118] = 16'd32597;
    assign memory[1119] = 16'd32594;
    assign memory[1120] = 16'd32590;
    assign memory[1121] = 16'd32586;
    assign memory[1122] = 16'd32583;
    assign memory[1123] = 16'd32579;
    assign memory[1124] = 16'd32575;
    assign memory[1125] = 16'd32571;
    assign memory[1126] = 16'd32567;
    assign memory[1127] = 16'd32563;
    assign memory[1128] = 16'd32559;
    assign memory[1129] = 16'd32555;
    assign memory[1130] = 16'd32551;
    assign memory[1131] = 16'd32547;
    assign memory[1132] = 16'd32543;
    assign memory[1133] = 16'd32539;
    assign memory[1134] = 16'd32535;
    assign memory[1135] = 16'd32531;
    assign memory[1136] = 16'd32526;
    assign memory[1137] = 16'd32522;
    assign memory[1138] = 16'd32518;
    assign memory[1139] = 16'd32513;
    assign memory[1140] = 16'd32509;
    assign memory[1141] = 16'd32504;
    assign memory[1142] = 16'd32500;
    assign memory[1143] = 16'd32495;
    assign memory[1144] = 16'd32491;
    assign memory[1145] = 16'd32486;
    assign memory[1146] = 16'd32481;
    assign memory[1147] = 16'd32477;
    assign memory[1148] = 16'd32472;
    assign memory[1149] = 16'd32467;
    assign memory[1150] = 16'd32462;
    assign memory[1151] = 16'd32458;
    assign memory[1152] = 16'd32453;
    assign memory[1153] = 16'd32448;
    assign memory[1154] = 16'd32443;
    assign memory[1155] = 16'd32438;
    assign memory[1156] = 16'd32433;
    assign memory[1157] = 16'd32428;
    assign memory[1158] = 16'd32423;
    assign memory[1159] = 16'd32417;
    assign memory[1160] = 16'd32412;
    assign memory[1161] = 16'd32407;
    assign memory[1162] = 16'd32402;
    assign memory[1163] = 16'd32396;
    assign memory[1164] = 16'd32391;
    assign memory[1165] = 16'd32386;
    assign memory[1166] = 16'd32380;
    assign memory[1167] = 16'd32375;
    assign memory[1168] = 16'd32369;
    assign memory[1169] = 16'd32364;
    assign memory[1170] = 16'd32358;
    assign memory[1171] = 16'd32353;
    assign memory[1172] = 16'd32347;
    assign memory[1173] = 16'd32341;
    assign memory[1174] = 16'd32336;
    assign memory[1175] = 16'd32330;
    assign memory[1176] = 16'd32324;
    assign memory[1177] = 16'd32318;
    assign memory[1178] = 16'd32312;
    assign memory[1179] = 16'd32307;
    assign memory[1180] = 16'd32301;
    assign memory[1181] = 16'd32295;
    assign memory[1182] = 16'd32289;
    assign memory[1183] = 16'd32283;
    assign memory[1184] = 16'd32276;
    assign memory[1185] = 16'd32270;
    assign memory[1186] = 16'd32264;
    assign memory[1187] = 16'd32258;
    assign memory[1188] = 16'd32252;
    assign memory[1189] = 16'd32245;
    assign memory[1190] = 16'd32239;
    assign memory[1191] = 16'd32233;
    assign memory[1192] = 16'd32226;
    assign memory[1193] = 16'd32220;
    assign memory[1194] = 16'd32214;
    assign memory[1195] = 16'd32207;
    assign memory[1196] = 16'd32201;
    assign memory[1197] = 16'd32194;
    assign memory[1198] = 16'd32187;
    assign memory[1199] = 16'd32181;
    assign memory[1200] = 16'd32174;
    assign memory[1201] = 16'd32167;
    assign memory[1202] = 16'd32161;
    assign memory[1203] = 16'd32154;
    assign memory[1204] = 16'd32147;
    assign memory[1205] = 16'd32140;
    assign memory[1206] = 16'd32133;
    assign memory[1207] = 16'd32126;
    assign memory[1208] = 16'd32119;
    assign memory[1209] = 16'd32112;
    assign memory[1210] = 16'd32105;
    assign memory[1211] = 16'd32098;
    assign memory[1212] = 16'd32091;
    assign memory[1213] = 16'd32084;
    assign memory[1214] = 16'd32077;
    assign memory[1215] = 16'd32069;
    assign memory[1216] = 16'd32062;
    assign memory[1217] = 16'd32055;
    assign memory[1218] = 16'd32047;
    assign memory[1219] = 16'd32040;
    assign memory[1220] = 16'd32033;
    assign memory[1221] = 16'd32025;
    assign memory[1222] = 16'd32018;
    assign memory[1223] = 16'd32010;
    assign memory[1224] = 16'd32002;
    assign memory[1225] = 16'd31995;
    assign memory[1226] = 16'd31987;
    assign memory[1227] = 16'd31980;
    assign memory[1228] = 16'd31972;
    assign memory[1229] = 16'd31964;
    assign memory[1230] = 16'd31956;
    assign memory[1231] = 16'd31948;
    assign memory[1232] = 16'd31941;
    assign memory[1233] = 16'd31933;
    assign memory[1234] = 16'd31925;
    assign memory[1235] = 16'd31917;
    assign memory[1236] = 16'd31909;
    assign memory[1237] = 16'd31901;
    assign memory[1238] = 16'd31893;
    assign memory[1239] = 16'd31884;
    assign memory[1240] = 16'd31876;
    assign memory[1241] = 16'd31868;
    assign memory[1242] = 16'd31860;
    assign memory[1243] = 16'd31852;
    assign memory[1244] = 16'd31843;
    assign memory[1245] = 16'd31835;
    assign memory[1246] = 16'd31827;
    assign memory[1247] = 16'd31818;
    assign memory[1248] = 16'd31810;
    assign memory[1249] = 16'd31801;
    assign memory[1250] = 16'd31793;
    assign memory[1251] = 16'd31784;
    assign memory[1252] = 16'd31776;
    assign memory[1253] = 16'd31767;
    assign memory[1254] = 16'd31758;
    assign memory[1255] = 16'd31750;
    assign memory[1256] = 16'd31741;
    assign memory[1257] = 16'd31732;
    assign memory[1258] = 16'd31723;
    assign memory[1259] = 16'd31714;
    assign memory[1260] = 16'd31706;
    assign memory[1261] = 16'd31697;
    assign memory[1262] = 16'd31688;
    assign memory[1263] = 16'd31679;
    assign memory[1264] = 16'd31670;
    assign memory[1265] = 16'd31661;
    assign memory[1266] = 16'd31651;
    assign memory[1267] = 16'd31642;
    assign memory[1268] = 16'd31633;
    assign memory[1269] = 16'd31624;
    assign memory[1270] = 16'd31615;
    assign memory[1271] = 16'd31605;
    assign memory[1272] = 16'd31596;
    assign memory[1273] = 16'd31587;
    assign memory[1274] = 16'd31577;
    assign memory[1275] = 16'd31568;
    assign memory[1276] = 16'd31559;
    assign memory[1277] = 16'd31549;
    assign memory[1278] = 16'd31540;
    assign memory[1279] = 16'd31530;
    assign memory[1280] = 16'd31520;
    assign memory[1281] = 16'd31511;
    assign memory[1282] = 16'd31501;
    assign memory[1283] = 16'd31491;
    assign memory[1284] = 16'd31482;
    assign memory[1285] = 16'd31472;
    assign memory[1286] = 16'd31462;
    assign memory[1287] = 16'd31452;
    assign memory[1288] = 16'd31442;
    assign memory[1289] = 16'd31432;
    assign memory[1290] = 16'd31422;
    assign memory[1291] = 16'd31412;
    assign memory[1292] = 16'd31402;
    assign memory[1293] = 16'd31392;
    assign memory[1294] = 16'd31382;
    assign memory[1295] = 16'd31372;
    assign memory[1296] = 16'd31362;
    assign memory[1297] = 16'd31352;
    assign memory[1298] = 16'd31341;
    assign memory[1299] = 16'd31331;
    assign memory[1300] = 16'd31321;
    assign memory[1301] = 16'd31311;
    assign memory[1302] = 16'd31300;
    assign memory[1303] = 16'd31290;
    assign memory[1304] = 16'd31279;
    assign memory[1305] = 16'd31269;
    assign memory[1306] = 16'd31258;
    assign memory[1307] = 16'd31248;
    assign memory[1308] = 16'd31237;
    assign memory[1309] = 16'd31227;
    assign memory[1310] = 16'd31216;
    assign memory[1311] = 16'd31205;
    assign memory[1312] = 16'd31194;
    assign memory[1313] = 16'd31184;
    assign memory[1314] = 16'd31173;
    assign memory[1315] = 16'd31162;
    assign memory[1316] = 16'd31151;
    assign memory[1317] = 16'd31140;
    assign memory[1318] = 16'd31129;
    assign memory[1319] = 16'd31118;
    assign memory[1320] = 16'd31107;
    assign memory[1321] = 16'd31096;
    assign memory[1322] = 16'd31085;
    assign memory[1323] = 16'd31074;
    assign memory[1324] = 16'd31063;
    assign memory[1325] = 16'd31052;
    assign memory[1326] = 16'd31041;
    assign memory[1327] = 16'd31029;
    assign memory[1328] = 16'd31018;
    assign memory[1329] = 16'd31007;
    assign memory[1330] = 16'd30995;
    assign memory[1331] = 16'd30984;
    assign memory[1332] = 16'd30973;
    assign memory[1333] = 16'd30961;
    assign memory[1334] = 16'd30950;
    assign memory[1335] = 16'd30938;
    assign memory[1336] = 16'd30927;
    assign memory[1337] = 16'd30915;
    assign memory[1338] = 16'd30903;
    assign memory[1339] = 16'd30892;
    assign memory[1340] = 16'd30880;
    assign memory[1341] = 16'd30868;
    assign memory[1342] = 16'd30857;
    assign memory[1343] = 16'd30845;
    assign memory[1344] = 16'd30833;
    assign memory[1345] = 16'd30821;
    assign memory[1346] = 16'd30809;
    assign memory[1347] = 16'd30797;
    assign memory[1348] = 16'd30785;
    assign memory[1349] = 16'd30773;
    assign memory[1350] = 16'd30761;
    assign memory[1351] = 16'd30749;
    assign memory[1352] = 16'd30737;
    assign memory[1353] = 16'd30725;
    assign memory[1354] = 16'd30713;
    assign memory[1355] = 16'd30701;
    assign memory[1356] = 16'd30688;
    assign memory[1357] = 16'd30676;
    assign memory[1358] = 16'd30664;
    assign memory[1359] = 16'd30651;
    assign memory[1360] = 16'd30639;
    assign memory[1361] = 16'd30627;
    assign memory[1362] = 16'd30614;
    assign memory[1363] = 16'd30602;
    assign memory[1364] = 16'd30589;
    assign memory[1365] = 16'd30577;
    assign memory[1366] = 16'd30564;
    assign memory[1367] = 16'd30551;
    assign memory[1368] = 16'd30539;
    assign memory[1369] = 16'd30526;
    assign memory[1370] = 16'd30513;
    assign memory[1371] = 16'd30501;
    assign memory[1372] = 16'd30488;
    assign memory[1373] = 16'd30475;
    assign memory[1374] = 16'd30462;
    assign memory[1375] = 16'd30449;
    assign memory[1376] = 16'd30437;
    assign memory[1377] = 16'd30424;
    assign memory[1378] = 16'd30411;
    assign memory[1379] = 16'd30398;
    assign memory[1380] = 16'd30385;
    assign memory[1381] = 16'd30372;
    assign memory[1382] = 16'd30358;
    assign memory[1383] = 16'd30345;
    assign memory[1384] = 16'd30332;
    assign memory[1385] = 16'd30319;
    assign memory[1386] = 16'd30306;
    assign memory[1387] = 16'd30292;
    assign memory[1388] = 16'd30279;
    assign memory[1389] = 16'd30266;
    assign memory[1390] = 16'd30252;
    assign memory[1391] = 16'd30239;
    assign memory[1392] = 16'd30226;
    assign memory[1393] = 16'd30212;
    assign memory[1394] = 16'd30199;
    assign memory[1395] = 16'd30185;
    assign memory[1396] = 16'd30172;
    assign memory[1397] = 16'd30158;
    assign memory[1398] = 16'd30144;
    assign memory[1399] = 16'd30131;
    assign memory[1400] = 16'd30117;
    assign memory[1401] = 16'd30103;
    assign memory[1402] = 16'd30089;
    assign memory[1403] = 16'd30076;
    assign memory[1404] = 16'd30062;
    assign memory[1405] = 16'd30048;
    assign memory[1406] = 16'd30034;
    assign memory[1407] = 16'd30020;
    assign memory[1408] = 16'd30006;
    assign memory[1409] = 16'd29992;
    assign memory[1410] = 16'd29978;
    assign memory[1411] = 16'd29964;
    assign memory[1412] = 16'd29950;
    assign memory[1413] = 16'd29936;
    assign memory[1414] = 16'd29922;
    assign memory[1415] = 16'd29908;
    assign memory[1416] = 16'd29894;
    assign memory[1417] = 16'd29879;
    assign memory[1418] = 16'd29865;
    assign memory[1419] = 16'd29851;
    assign memory[1420] = 16'd29836;
    assign memory[1421] = 16'd29822;
    assign memory[1422] = 16'd29808;
    assign memory[1423] = 16'd29793;
    assign memory[1424] = 16'd29779;
    assign memory[1425] = 16'd29764;
    assign memory[1426] = 16'd29750;
    assign memory[1427] = 16'd29735;
    assign memory[1428] = 16'd29721;
    assign memory[1429] = 16'd29706;
    assign memory[1430] = 16'd29691;
    assign memory[1431] = 16'd29677;
    assign memory[1432] = 16'd29662;
    assign memory[1433] = 16'd29647;
    assign memory[1434] = 16'd29633;
    assign memory[1435] = 16'd29618;
    assign memory[1436] = 16'd29603;
    assign memory[1437] = 16'd29588;
    assign memory[1438] = 16'd29573;
    assign memory[1439] = 16'd29558;
    assign memory[1440] = 16'd29543;
    assign memory[1441] = 16'd29528;
    assign memory[1442] = 16'd29513;
    assign memory[1443] = 16'd29498;
    assign memory[1444] = 16'd29483;
    assign memory[1445] = 16'd29468;
    assign memory[1446] = 16'd29453;
    assign memory[1447] = 16'd29438;
    assign memory[1448] = 16'd29422;
    assign memory[1449] = 16'd29407;
    assign memory[1450] = 16'd29392;
    assign memory[1451] = 16'd29377;
    assign memory[1452] = 16'd29361;
    assign memory[1453] = 16'd29346;
    assign memory[1454] = 16'd29331;
    assign memory[1455] = 16'd29315;
    assign memory[1456] = 16'd29300;
    assign memory[1457] = 16'd29284;
    assign memory[1458] = 16'd29269;
    assign memory[1459] = 16'd29253;
    assign memory[1460] = 16'd29238;
    assign memory[1461] = 16'd29222;
    assign memory[1462] = 16'd29206;
    assign memory[1463] = 16'd29191;
    assign memory[1464] = 16'd29175;
    assign memory[1465] = 16'd29159;
    assign memory[1466] = 16'd29144;
    assign memory[1467] = 16'd29128;
    assign memory[1468] = 16'd29112;
    assign memory[1469] = 16'd29096;
    assign memory[1470] = 16'd29080;
    assign memory[1471] = 16'd29064;
    assign memory[1472] = 16'd29049;
    assign memory[1473] = 16'd29033;
    assign memory[1474] = 16'd29017;
    assign memory[1475] = 16'd29001;
    assign memory[1476] = 16'd28984;
    assign memory[1477] = 16'd28968;
    assign memory[1478] = 16'd28952;
    assign memory[1479] = 16'd28936;
    assign memory[1480] = 16'd28920;
    assign memory[1481] = 16'd28904;
    assign memory[1482] = 16'd28888;
    assign memory[1483] = 16'd28871;
    assign memory[1484] = 16'd28855;
    assign memory[1485] = 16'd28839;
    assign memory[1486] = 16'd28822;
    assign memory[1487] = 16'd28806;
    assign memory[1488] = 16'd28790;
    assign memory[1489] = 16'd28773;
    assign memory[1490] = 16'd28757;
    assign memory[1491] = 16'd28740;
    assign memory[1492] = 16'd28724;
    assign memory[1493] = 16'd28707;
    assign memory[1494] = 16'd28691;
    assign memory[1495] = 16'd28674;
    assign memory[1496] = 16'd28657;
    assign memory[1497] = 16'd28641;
    assign memory[1498] = 16'd28624;
    assign memory[1499] = 16'd28607;
    assign memory[1500] = 16'd28591;
    assign memory[1501] = 16'd28574;
    assign memory[1502] = 16'd28557;
    assign memory[1503] = 16'd28540;
    assign memory[1504] = 16'd28523;
    assign memory[1505] = 16'd28506;
    assign memory[1506] = 16'd28489;
    assign memory[1507] = 16'd28472;
    assign memory[1508] = 16'd28456;
    assign memory[1509] = 16'd28438;
    assign memory[1510] = 16'd28421;
    assign memory[1511] = 16'd28404;
    assign memory[1512] = 16'd28387;
    assign memory[1513] = 16'd28370;
    assign memory[1514] = 16'd28353;
    assign memory[1515] = 16'd28336;
    assign memory[1516] = 16'd28319;
    assign memory[1517] = 16'd28301;
    assign memory[1518] = 16'd28284;
    assign memory[1519] = 16'd28267;
    assign memory[1520] = 16'd28250;
    assign memory[1521] = 16'd28232;
    assign memory[1522] = 16'd28215;
    assign memory[1523] = 16'd28197;
    assign memory[1524] = 16'd28180;
    assign memory[1525] = 16'd28163;
    assign memory[1526] = 16'd28145;
    assign memory[1527] = 16'd28128;
    assign memory[1528] = 16'd28110;
    assign memory[1529] = 16'd28092;
    assign memory[1530] = 16'd28075;
    assign memory[1531] = 16'd28057;
    assign memory[1532] = 16'd28040;
    assign memory[1533] = 16'd28022;
    assign memory[1534] = 16'd28004;
    assign memory[1535] = 16'd27986;
    assign memory[1536] = 16'd27969;
    assign memory[1537] = 16'd27951;
    assign memory[1538] = 16'd27933;
    assign memory[1539] = 16'd27915;
    assign memory[1540] = 16'd27897;
    assign memory[1541] = 16'd27880;
    assign memory[1542] = 16'd27862;
    assign memory[1543] = 16'd27844;
    assign memory[1544] = 16'd27826;
    assign memory[1545] = 16'd27808;
    assign memory[1546] = 16'd27790;
    assign memory[1547] = 16'd27772;
    assign memory[1548] = 16'd27754;
    assign memory[1549] = 16'd27735;
    assign memory[1550] = 16'd27717;
    assign memory[1551] = 16'd27699;
    assign memory[1552] = 16'd27681;
    assign memory[1553] = 16'd27663;
    assign memory[1554] = 16'd27644;
    assign memory[1555] = 16'd27626;
    assign memory[1556] = 16'd27608;
    assign memory[1557] = 16'd27590;
    assign memory[1558] = 16'd27571;
    assign memory[1559] = 16'd27553;
    assign memory[1560] = 16'd27534;
    assign memory[1561] = 16'd27516;
    assign memory[1562] = 16'd27498;
    assign memory[1563] = 16'd27479;
    assign memory[1564] = 16'd27461;
    assign memory[1565] = 16'd27442;
    assign memory[1566] = 16'd27424;
    assign memory[1567] = 16'd27405;
    assign memory[1568] = 16'd27386;
    assign memory[1569] = 16'd27368;
    assign memory[1570] = 16'd27349;
    assign memory[1571] = 16'd27330;
    assign memory[1572] = 16'd27312;
    assign memory[1573] = 16'd27293;
    assign memory[1574] = 16'd27274;
    assign memory[1575] = 16'd27255;
    assign memory[1576] = 16'd27237;
    assign memory[1577] = 16'd27218;
    assign memory[1578] = 16'd27199;
    assign memory[1579] = 16'd27180;
    assign memory[1580] = 16'd27161;
    assign memory[1581] = 16'd27142;
    assign memory[1582] = 16'd27123;
    assign memory[1583] = 16'd27104;
    assign memory[1584] = 16'd27085;
    assign memory[1585] = 16'd27066;
    assign memory[1586] = 16'd27047;
    assign memory[1587] = 16'd27028;
    assign memory[1588] = 16'd27009;
    assign memory[1589] = 16'd26990;
    assign memory[1590] = 16'd26970;
    assign memory[1591] = 16'd26951;
    assign memory[1592] = 16'd26932;
    assign memory[1593] = 16'd26913;
    assign memory[1594] = 16'd26894;
    assign memory[1595] = 16'd26874;
    assign memory[1596] = 16'd26855;
    assign memory[1597] = 16'd26836;
    assign memory[1598] = 16'd26816;
    assign memory[1599] = 16'd26797;
    assign memory[1600] = 16'd26777;
    assign memory[1601] = 16'd26758;
    assign memory[1602] = 16'd26738;
    assign memory[1603] = 16'd26719;
    assign memory[1604] = 16'd26699;
    assign memory[1605] = 16'd26680;
    assign memory[1606] = 16'd26660;
    assign memory[1607] = 16'd26641;
    assign memory[1608] = 16'd26621;
    assign memory[1609] = 16'd26602;
    assign memory[1610] = 16'd26582;
    assign memory[1611] = 16'd26562;
    assign memory[1612] = 16'd26543;
    assign memory[1613] = 16'd26523;
    assign memory[1614] = 16'd26503;
    assign memory[1615] = 16'd26483;
    assign memory[1616] = 16'd26463;
    assign memory[1617] = 16'd26444;
    assign memory[1618] = 16'd26424;
    assign memory[1619] = 16'd26404;
    assign memory[1620] = 16'd26384;
    assign memory[1621] = 16'd26364;
    assign memory[1622] = 16'd26344;
    assign memory[1623] = 16'd26324;
    assign memory[1624] = 16'd26304;
    assign memory[1625] = 16'd26284;
    assign memory[1626] = 16'd26264;
    assign memory[1627] = 16'd26244;
    assign memory[1628] = 16'd26224;
    assign memory[1629] = 16'd26204;
    assign memory[1630] = 16'd26184;
    assign memory[1631] = 16'd26164;
    assign memory[1632] = 16'd26143;
    assign memory[1633] = 16'd26123;
    assign memory[1634] = 16'd26103;
    assign memory[1635] = 16'd26083;
    assign memory[1636] = 16'd26063;
    assign memory[1637] = 16'd26042;
    assign memory[1638] = 16'd26022;
    assign memory[1639] = 16'd26002;
    assign memory[1640] = 16'd25981;
    assign memory[1641] = 16'd25961;
    assign memory[1642] = 16'd25940;
    assign memory[1643] = 16'd25920;
    assign memory[1644] = 16'd25900;
    assign memory[1645] = 16'd25879;
    assign memory[1646] = 16'd25859;
    assign memory[1647] = 16'd25838;
    assign memory[1648] = 16'd25818;
    assign memory[1649] = 16'd25797;
    assign memory[1650] = 16'd25776;
    assign memory[1651] = 16'd25756;
    assign memory[1652] = 16'd25735;
    assign memory[1653] = 16'd25715;
    assign memory[1654] = 16'd25694;
    assign memory[1655] = 16'd25673;
    assign memory[1656] = 16'd25652;
    assign memory[1657] = 16'd25632;
    assign memory[1658] = 16'd25611;
    assign memory[1659] = 16'd25590;
    assign memory[1660] = 16'd25569;
    assign memory[1661] = 16'd25549;
    assign memory[1662] = 16'd25528;
    assign memory[1663] = 16'd25507;
    assign memory[1664] = 16'd25486;
    assign memory[1665] = 16'd25465;
    assign memory[1666] = 16'd25444;
    assign memory[1667] = 16'd25423;
    assign memory[1668] = 16'd25402;
    assign memory[1669] = 16'd25381;
    assign memory[1670] = 16'd25360;
    assign memory[1671] = 16'd25339;
    assign memory[1672] = 16'd25318;
    assign memory[1673] = 16'd25297;
    assign memory[1674] = 16'd25276;
    assign memory[1675] = 16'd25255;
    assign memory[1676] = 16'd25234;
    assign memory[1677] = 16'd25213;
    assign memory[1678] = 16'd25191;
    assign memory[1679] = 16'd25170;
    assign memory[1680] = 16'd25149;
    assign memory[1681] = 16'd25128;
    assign memory[1682] = 16'd25106;
    assign memory[1683] = 16'd25085;
    assign memory[1684] = 16'd25064;
    assign memory[1685] = 16'd25042;
    assign memory[1686] = 16'd25021;
    assign memory[1687] = 16'd25000;
    assign memory[1688] = 16'd24978;
    assign memory[1689] = 16'd24957;
    assign memory[1690] = 16'd24936;
    assign memory[1691] = 16'd24914;
    assign memory[1692] = 16'd24893;
    assign memory[1693] = 16'd24871;
    assign memory[1694] = 16'd24850;
    assign memory[1695] = 16'd24828;
    assign memory[1696] = 16'd24807;
    assign memory[1697] = 16'd24785;
    assign memory[1698] = 16'd24763;
    assign memory[1699] = 16'd24742;
    assign memory[1700] = 16'd24720;
    assign memory[1701] = 16'd24699;
    assign memory[1702] = 16'd24677;
    assign memory[1703] = 16'd24655;
    assign memory[1704] = 16'd24633;
    assign memory[1705] = 16'd24612;
    assign memory[1706] = 16'd24590;
    assign memory[1707] = 16'd24568;
    assign memory[1708] = 16'd24546;
    assign memory[1709] = 16'd24525;
    assign memory[1710] = 16'd24503;
    assign memory[1711] = 16'd24481;
    assign memory[1712] = 16'd24459;
    assign memory[1713] = 16'd24437;
    assign memory[1714] = 16'd24415;
    assign memory[1715] = 16'd24393;
    assign memory[1716] = 16'd24372;
    assign memory[1717] = 16'd24350;
    assign memory[1718] = 16'd24328;
    assign memory[1719] = 16'd24306;
    assign memory[1720] = 16'd24284;
    assign memory[1721] = 16'd24262;
    assign memory[1722] = 16'd24240;
    assign memory[1723] = 16'd24217;
    assign memory[1724] = 16'd24195;
    assign memory[1725] = 16'd24173;
    assign memory[1726] = 16'd24151;
    assign memory[1727] = 16'd24129;
    assign memory[1728] = 16'd24107;
    assign memory[1729] = 16'd24085;
    assign memory[1730] = 16'd24062;
    assign memory[1731] = 16'd24040;
    assign memory[1732] = 16'd24018;
    assign memory[1733] = 16'd23996;
    assign memory[1734] = 16'd23974;
    assign memory[1735] = 16'd23951;
    assign memory[1736] = 16'd23929;
    assign memory[1737] = 16'd23907;
    assign memory[1738] = 16'd23884;
    assign memory[1739] = 16'd23862;
    assign memory[1740] = 16'd23840;
    assign memory[1741] = 16'd23817;
    assign memory[1742] = 16'd23795;
    assign memory[1743] = 16'd23772;
    assign memory[1744] = 16'd23750;
    assign memory[1745] = 16'd23727;
    assign memory[1746] = 16'd23705;
    assign memory[1747] = 16'd23683;
    assign memory[1748] = 16'd23660;
    assign memory[1749] = 16'd23637;
    assign memory[1750] = 16'd23615;
    assign memory[1751] = 16'd23592;
    assign memory[1752] = 16'd23570;
    assign memory[1753] = 16'd23547;
    assign memory[1754] = 16'd23525;
    assign memory[1755] = 16'd23502;
    assign memory[1756] = 16'd23479;
    assign memory[1757] = 16'd23457;
    assign memory[1758] = 16'd23434;
    assign memory[1759] = 16'd23411;
    assign memory[1760] = 16'd23389;
    assign memory[1761] = 16'd23366;
    assign memory[1762] = 16'd23343;
    assign memory[1763] = 16'd23320;
    assign memory[1764] = 16'd23298;
    assign memory[1765] = 16'd23275;
    assign memory[1766] = 16'd23252;
    assign memory[1767] = 16'd23229;
    assign memory[1768] = 16'd23206;
    assign memory[1769] = 16'd23183;
    assign memory[1770] = 16'd23161;
    assign memory[1771] = 16'd23138;
    assign memory[1772] = 16'd23115;
    assign memory[1773] = 16'd23092;
    assign memory[1774] = 16'd23069;
    assign memory[1775] = 16'd23046;
    assign memory[1776] = 16'd23023;
    assign memory[1777] = 16'd23000;
    assign memory[1778] = 16'd22977;
    assign memory[1779] = 16'd22954;
    assign memory[1780] = 16'd22931;
    assign memory[1781] = 16'd22908;
    assign memory[1782] = 16'd22885;
    assign memory[1783] = 16'd22862;
    assign memory[1784] = 16'd22839;
    assign memory[1785] = 16'd22816;
    assign memory[1786] = 16'd22792;
    assign memory[1787] = 16'd22769;
    assign memory[1788] = 16'd22746;
    assign memory[1789] = 16'd22723;
    assign memory[1790] = 16'd22700;
    assign memory[1791] = 16'd22677;
    assign memory[1792] = 16'd22653;
    assign memory[1793] = 16'd22630;
    assign memory[1794] = 16'd22607;
    assign memory[1795] = 16'd22584;
    assign memory[1796] = 16'd22560;
    assign memory[1797] = 16'd22537;
    assign memory[1798] = 16'd22514;
    assign memory[1799] = 16'd22490;
    assign memory[1800] = 16'd22467;
    assign memory[1801] = 16'd22444;
    assign memory[1802] = 16'd22420;
    assign memory[1803] = 16'd22397;
    assign memory[1804] = 16'd22374;
    assign memory[1805] = 16'd22350;
    assign memory[1806] = 16'd22327;
    assign memory[1807] = 16'd22303;
    assign memory[1808] = 16'd22280;
    assign memory[1809] = 16'd22257;
    assign memory[1810] = 16'd22233;
    assign memory[1811] = 16'd22210;
    assign memory[1812] = 16'd22186;
    assign memory[1813] = 16'd22163;
    assign memory[1814] = 16'd22139;
    assign memory[1815] = 16'd22116;
    assign memory[1816] = 16'd22092;
    assign memory[1817] = 16'd22068;
    assign memory[1818] = 16'd22045;
    assign memory[1819] = 16'd22021;
    assign memory[1820] = 16'd21998;
    assign memory[1821] = 16'd21974;
    assign memory[1822] = 16'd21950;
    assign memory[1823] = 16'd21927;
    assign memory[1824] = 16'd21903;
    assign memory[1825] = 16'd21879;
    assign memory[1826] = 16'd21856;
    assign memory[1827] = 16'd21832;
    assign memory[1828] = 16'd21808;
    assign memory[1829] = 16'd21785;
    assign memory[1830] = 16'd21761;
    assign memory[1831] = 16'd21737;
    assign memory[1832] = 16'd21713;
    assign memory[1833] = 16'd21690;
    assign memory[1834] = 16'd21666;
    assign memory[1835] = 16'd21642;
    assign memory[1836] = 16'd21618;
    assign memory[1837] = 16'd21594;
    assign memory[1838] = 16'd21571;
    assign memory[1839] = 16'd21547;
    assign memory[1840] = 16'd21523;
    assign memory[1841] = 16'd21499;
    assign memory[1842] = 16'd21475;
    assign memory[1843] = 16'd21451;
    assign memory[1844] = 16'd21427;
    assign memory[1845] = 16'd21403;
    assign memory[1846] = 16'd21379;
    assign memory[1847] = 16'd21356;
    assign memory[1848] = 16'd21332;
    assign memory[1849] = 16'd21308;
    assign memory[1850] = 16'd21284;
    assign memory[1851] = 16'd21260;
    assign memory[1852] = 16'd21236;
    assign memory[1853] = 16'd21212;
    assign memory[1854] = 16'd21188;
    assign memory[1855] = 16'd21164;
    assign memory[1856] = 16'd21140;
    assign memory[1857] = 16'd21115;
    assign memory[1858] = 16'd21091;
    assign memory[1859] = 16'd21067;
    assign memory[1860] = 16'd21043;
    assign memory[1861] = 16'd21019;
    assign memory[1862] = 16'd20995;
    assign memory[1863] = 16'd20971;
    assign memory[1864] = 16'd20947;
    assign memory[1865] = 16'd20923;
    assign memory[1866] = 16'd20898;
    assign memory[1867] = 16'd20874;
    assign memory[1868] = 16'd20850;
    assign memory[1869] = 16'd20826;
    assign memory[1870] = 16'd20802;
    assign memory[1871] = 16'd20778;
    assign memory[1872] = 16'd20753;
    assign memory[1873] = 16'd20729;
    assign memory[1874] = 16'd20705;
    assign memory[1875] = 16'd20681;
    assign memory[1876] = 16'd20656;
    assign memory[1877] = 16'd20632;
    assign memory[1878] = 16'd20608;
    assign memory[1879] = 16'd20584;
    assign memory[1880] = 16'd20559;
    assign memory[1881] = 16'd20535;
    assign memory[1882] = 16'd20511;
    assign memory[1883] = 16'd20486;
    assign memory[1884] = 16'd20462;
    assign memory[1885] = 16'd20438;
    assign memory[1886] = 16'd20413;
    assign memory[1887] = 16'd20389;
    assign memory[1888] = 16'd20364;
    assign memory[1889] = 16'd20340;
    assign memory[1890] = 16'd20316;
    assign memory[1891] = 16'd20291;
    assign memory[1892] = 16'd20267;
    assign memory[1893] = 16'd20242;
    assign memory[1894] = 16'd20218;
    assign memory[1895] = 16'd20194;
    assign memory[1896] = 16'd20169;
    assign memory[1897] = 16'd20145;
    assign memory[1898] = 16'd20120;
    assign memory[1899] = 16'd20096;
    assign memory[1900] = 16'd20071;
    assign memory[1901] = 16'd20047;
    assign memory[1902] = 16'd20022;
    assign memory[1903] = 16'd19998;
    assign memory[1904] = 16'd19973;
    assign memory[1905] = 16'd19949;
    assign memory[1906] = 16'd19924;
    assign memory[1907] = 16'd19900;
    assign memory[1908] = 16'd19875;
    assign memory[1909] = 16'd19851;
    assign memory[1910] = 16'd19826;
    assign memory[1911] = 16'd19801;
    assign memory[1912] = 16'd19777;
    assign memory[1913] = 16'd19752;
    assign memory[1914] = 16'd19728;
    assign memory[1915] = 16'd19703;
    assign memory[1916] = 16'd19678;
    assign memory[1917] = 16'd19654;
    assign memory[1918] = 16'd19629;
    assign memory[1919] = 16'd19605;
    assign memory[1920] = 16'd19580;
    assign memory[1921] = 16'd19555;
    assign memory[1922] = 16'd19531;
    assign memory[1923] = 16'd19506;
    assign memory[1924] = 16'd19481;
    assign memory[1925] = 16'd19457;
    assign memory[1926] = 16'd19432;
    assign memory[1927] = 16'd19407;
    assign memory[1928] = 16'd19382;
    assign memory[1929] = 16'd19358;
    assign memory[1930] = 16'd19333;
    assign memory[1931] = 16'd19308;
    assign memory[1932] = 16'd19284;
    assign memory[1933] = 16'd19259;
    assign memory[1934] = 16'd19234;
    assign memory[1935] = 16'd19209;
    assign memory[1936] = 16'd19185;
    assign memory[1937] = 16'd19160;
    assign memory[1938] = 16'd19135;
    assign memory[1939] = 16'd19110;
    assign memory[1940] = 16'd19085;
    assign memory[1941] = 16'd19061;
    assign memory[1942] = 16'd19036;
    assign memory[1943] = 16'd19011;
    assign memory[1944] = 16'd18986;
    assign memory[1945] = 16'd18961;
    assign memory[1946] = 16'd18937;
    assign memory[1947] = 16'd18912;
    assign memory[1948] = 16'd18887;
    assign memory[1949] = 16'd18862;
    assign memory[1950] = 16'd18837;
    assign memory[1951] = 16'd18812;
    assign memory[1952] = 16'd18788;
    assign memory[1953] = 16'd18763;
    assign memory[1954] = 16'd18738;
    assign memory[1955] = 16'd18713;
    assign memory[1956] = 16'd18688;
    assign memory[1957] = 16'd18663;
    assign memory[1958] = 16'd18638;
    assign memory[1959] = 16'd18613;
    assign memory[1960] = 16'd18588;
    assign memory[1961] = 16'd18564;
    assign memory[1962] = 16'd18539;
    assign memory[1963] = 16'd18514;
    assign memory[1964] = 16'd18489;
    assign memory[1965] = 16'd18464;
    assign memory[1966] = 16'd18439;
    assign memory[1967] = 16'd18414;
    assign memory[1968] = 16'd18389;
    assign memory[1969] = 16'd18364;
    assign memory[1970] = 16'd18339;
    assign memory[1971] = 16'd18314;
    assign memory[1972] = 16'd18289;
    assign memory[1973] = 16'd18264;
    assign memory[1974] = 16'd18239;
    assign memory[1975] = 16'd18214;
    assign memory[1976] = 16'd18189;
    assign memory[1977] = 16'd18164;
    assign memory[1978] = 16'd18139;
    assign memory[1979] = 16'd18114;
    assign memory[1980] = 16'd18089;
    assign memory[1981] = 16'd18064;
    assign memory[1982] = 16'd18039;
    assign memory[1983] = 16'd18014;
    assign memory[1984] = 16'd17989;
    assign memory[1985] = 16'd17964;
    assign memory[1986] = 16'd17939;
    assign memory[1987] = 16'd17914;
    assign memory[1988] = 16'd17889;
    assign memory[1989] = 16'd17864;
    assign memory[1990] = 16'd17839;
    assign memory[1991] = 16'd17814;
    assign memory[1992] = 16'd17789;
    assign memory[1993] = 16'd17764;
    assign memory[1994] = 16'd17739;
    assign memory[1995] = 16'd17714;
    assign memory[1996] = 16'd17689;
    assign memory[1997] = 16'd17664;
    assign memory[1998] = 16'd17639;
    assign memory[1999] = 16'd17614;
    assign memory[2000] = 16'd17589;
    assign memory[2001] = 16'd17564;
    assign memory[2002] = 16'd17539;
    assign memory[2003] = 16'd17514;
    assign memory[2004] = 16'd17489;
    assign memory[2005] = 16'd17463;
    assign memory[2006] = 16'd17438;
    assign memory[2007] = 16'd17413;
    assign memory[2008] = 16'd17388;
    assign memory[2009] = 16'd17363;
    assign memory[2010] = 16'd17338;
    assign memory[2011] = 16'd17313;
    assign memory[2012] = 16'd17288;
    assign memory[2013] = 16'd17263;
    assign memory[2014] = 16'd17238;
    assign memory[2015] = 16'd17213;
    assign memory[2016] = 16'd17187;
    assign memory[2017] = 16'd17162;
    assign memory[2018] = 16'd17137;
    assign memory[2019] = 16'd17112;
    assign memory[2020] = 16'd17087;
    assign memory[2021] = 16'd17062;
    assign memory[2022] = 16'd17037;
    assign memory[2023] = 16'd17012;
    assign memory[2024] = 16'd16987;
    assign memory[2025] = 16'd16961;
    assign memory[2026] = 16'd16936;
    assign memory[2027] = 16'd16911;
    assign memory[2028] = 16'd16886;
    assign memory[2029] = 16'd16861;
    assign memory[2030] = 16'd16836;
    assign memory[2031] = 16'd16811;
    assign memory[2032] = 16'd16786;
    assign memory[2033] = 16'd16760;
    assign memory[2034] = 16'd16735;
    assign memory[2035] = 16'd16710;
    assign memory[2036] = 16'd16685;
    assign memory[2037] = 16'd16660;
    assign memory[2038] = 16'd16635;
    assign memory[2039] = 16'd16610;
    assign memory[2040] = 16'd16585;
    assign memory[2041] = 16'd16559;
    assign memory[2042] = 16'd16534;
    assign memory[2043] = 16'd16509;
    assign memory[2044] = 16'd16484;
    assign memory[2045] = 16'd16459;
    assign memory[2046] = 16'd16434;
    assign memory[2047] = 16'd16409;
    assign memory[2048] = 16'd16384;
    assign memory[2049] = 16'd16359;
    assign memory[2050] = 16'd16334;
    assign memory[2051] = 16'd16309;
    assign memory[2052] = 16'd16284;
    assign memory[2053] = 16'd16259;
    assign memory[2054] = 16'd16234;
    assign memory[2055] = 16'd16209;
    assign memory[2056] = 16'd16183;
    assign memory[2057] = 16'd16158;
    assign memory[2058] = 16'd16133;
    assign memory[2059] = 16'd16108;
    assign memory[2060] = 16'd16083;
    assign memory[2061] = 16'd16058;
    assign memory[2062] = 16'd16033;
    assign memory[2063] = 16'd16008;
    assign memory[2064] = 16'd15982;
    assign memory[2065] = 16'd15957;
    assign memory[2066] = 16'd15932;
    assign memory[2067] = 16'd15907;
    assign memory[2068] = 16'd15882;
    assign memory[2069] = 16'd15857;
    assign memory[2070] = 16'd15832;
    assign memory[2071] = 16'd15807;
    assign memory[2072] = 16'd15781;
    assign memory[2073] = 16'd15756;
    assign memory[2074] = 16'd15731;
    assign memory[2075] = 16'd15706;
    assign memory[2076] = 16'd15681;
    assign memory[2077] = 16'd15656;
    assign memory[2078] = 16'd15631;
    assign memory[2079] = 16'd15606;
    assign memory[2080] = 16'd15581;
    assign memory[2081] = 16'd15555;
    assign memory[2082] = 16'd15530;
    assign memory[2083] = 16'd15505;
    assign memory[2084] = 16'd15480;
    assign memory[2085] = 16'd15455;
    assign memory[2086] = 16'd15430;
    assign memory[2087] = 16'd15405;
    assign memory[2088] = 16'd15380;
    assign memory[2089] = 16'd15355;
    assign memory[2090] = 16'd15330;
    assign memory[2091] = 16'd15305;
    assign memory[2092] = 16'd15279;
    assign memory[2093] = 16'd15254;
    assign memory[2094] = 16'd15229;
    assign memory[2095] = 16'd15204;
    assign memory[2096] = 16'd15179;
    assign memory[2097] = 16'd15154;
    assign memory[2098] = 16'd15129;
    assign memory[2099] = 16'd15104;
    assign memory[2100] = 16'd15079;
    assign memory[2101] = 16'd15054;
    assign memory[2102] = 16'd15029;
    assign memory[2103] = 16'd15004;
    assign memory[2104] = 16'd14979;
    assign memory[2105] = 16'd14954;
    assign memory[2106] = 16'd14929;
    assign memory[2107] = 16'd14904;
    assign memory[2108] = 16'd14879;
    assign memory[2109] = 16'd14854;
    assign memory[2110] = 16'd14829;
    assign memory[2111] = 16'd14804;
    assign memory[2112] = 16'd14779;
    assign memory[2113] = 16'd14754;
    assign memory[2114] = 16'd14729;
    assign memory[2115] = 16'd14704;
    assign memory[2116] = 16'd14679;
    assign memory[2117] = 16'd14654;
    assign memory[2118] = 16'd14629;
    assign memory[2119] = 16'd14604;
    assign memory[2120] = 16'd14579;
    assign memory[2121] = 16'd14554;
    assign memory[2122] = 16'd14529;
    assign memory[2123] = 16'd14504;
    assign memory[2124] = 16'd14479;
    assign memory[2125] = 16'd14454;
    assign memory[2126] = 16'd14429;
    assign memory[2127] = 16'd14404;
    assign memory[2128] = 16'd14379;
    assign memory[2129] = 16'd14354;
    assign memory[2130] = 16'd14329;
    assign memory[2131] = 16'd14304;
    assign memory[2132] = 16'd14279;
    assign memory[2133] = 16'd14254;
    assign memory[2134] = 16'd14229;
    assign memory[2135] = 16'd14204;
    assign memory[2136] = 16'd14180;
    assign memory[2137] = 16'd14155;
    assign memory[2138] = 16'd14130;
    assign memory[2139] = 16'd14105;
    assign memory[2140] = 16'd14080;
    assign memory[2141] = 16'd14055;
    assign memory[2142] = 16'd14030;
    assign memory[2143] = 16'd14005;
    assign memory[2144] = 16'd13980;
    assign memory[2145] = 16'd13956;
    assign memory[2146] = 16'd13931;
    assign memory[2147] = 16'd13906;
    assign memory[2148] = 16'd13881;
    assign memory[2149] = 16'd13856;
    assign memory[2150] = 16'd13831;
    assign memory[2151] = 16'd13807;
    assign memory[2152] = 16'd13782;
    assign memory[2153] = 16'd13757;
    assign memory[2154] = 16'd13732;
    assign memory[2155] = 16'd13707;
    assign memory[2156] = 16'd13683;
    assign memory[2157] = 16'd13658;
    assign memory[2158] = 16'd13633;
    assign memory[2159] = 16'd13608;
    assign memory[2160] = 16'd13583;
    assign memory[2161] = 16'd13559;
    assign memory[2162] = 16'd13534;
    assign memory[2163] = 16'd13509;
    assign memory[2164] = 16'd13484;
    assign memory[2165] = 16'd13460;
    assign memory[2166] = 16'd13435;
    assign memory[2167] = 16'd13410;
    assign memory[2168] = 16'd13386;
    assign memory[2169] = 16'd13361;
    assign memory[2170] = 16'd13336;
    assign memory[2171] = 16'd13311;
    assign memory[2172] = 16'd13287;
    assign memory[2173] = 16'd13262;
    assign memory[2174] = 16'd13237;
    assign memory[2175] = 16'd13213;
    assign memory[2176] = 16'd13188;
    assign memory[2177] = 16'd13163;
    assign memory[2178] = 16'd13139;
    assign memory[2179] = 16'd13114;
    assign memory[2180] = 16'd13090;
    assign memory[2181] = 16'd13065;
    assign memory[2182] = 16'd13040;
    assign memory[2183] = 16'd13016;
    assign memory[2184] = 16'd12991;
    assign memory[2185] = 16'd12967;
    assign memory[2186] = 16'd12942;
    assign memory[2187] = 16'd12917;
    assign memory[2188] = 16'd12893;
    assign memory[2189] = 16'd12868;
    assign memory[2190] = 16'd12844;
    assign memory[2191] = 16'd12819;
    assign memory[2192] = 16'd12795;
    assign memory[2193] = 16'd12770;
    assign memory[2194] = 16'd12746;
    assign memory[2195] = 16'd12721;
    assign memory[2196] = 16'd12697;
    assign memory[2197] = 16'd12672;
    assign memory[2198] = 16'd12648;
    assign memory[2199] = 16'd12623;
    assign memory[2200] = 16'd12599;
    assign memory[2201] = 16'd12574;
    assign memory[2202] = 16'd12550;
    assign memory[2203] = 16'd12526;
    assign memory[2204] = 16'd12501;
    assign memory[2205] = 16'd12477;
    assign memory[2206] = 16'd12452;
    assign memory[2207] = 16'd12428;
    assign memory[2208] = 16'd12404;
    assign memory[2209] = 16'd12379;
    assign memory[2210] = 16'd12355;
    assign memory[2211] = 16'd12330;
    assign memory[2212] = 16'd12306;
    assign memory[2213] = 16'd12282;
    assign memory[2214] = 16'd12257;
    assign memory[2215] = 16'd12233;
    assign memory[2216] = 16'd12209;
    assign memory[2217] = 16'd12184;
    assign memory[2218] = 16'd12160;
    assign memory[2219] = 16'd12136;
    assign memory[2220] = 16'd12112;
    assign memory[2221] = 16'd12087;
    assign memory[2222] = 16'd12063;
    assign memory[2223] = 16'd12039;
    assign memory[2224] = 16'd12015;
    assign memory[2225] = 16'd11990;
    assign memory[2226] = 16'd11966;
    assign memory[2227] = 16'd11942;
    assign memory[2228] = 16'd11918;
    assign memory[2229] = 16'd11894;
    assign memory[2230] = 16'd11870;
    assign memory[2231] = 16'd11845;
    assign memory[2232] = 16'd11821;
    assign memory[2233] = 16'd11797;
    assign memory[2234] = 16'd11773;
    assign memory[2235] = 16'd11749;
    assign memory[2236] = 16'd11725;
    assign memory[2237] = 16'd11701;
    assign memory[2238] = 16'd11677;
    assign memory[2239] = 16'd11653;
    assign memory[2240] = 16'd11628;
    assign memory[2241] = 16'd11604;
    assign memory[2242] = 16'd11580;
    assign memory[2243] = 16'd11556;
    assign memory[2244] = 16'd11532;
    assign memory[2245] = 16'd11508;
    assign memory[2246] = 16'd11484;
    assign memory[2247] = 16'd11460;
    assign memory[2248] = 16'd11436;
    assign memory[2249] = 16'd11412;
    assign memory[2250] = 16'd11389;
    assign memory[2251] = 16'd11365;
    assign memory[2252] = 16'd11341;
    assign memory[2253] = 16'd11317;
    assign memory[2254] = 16'd11293;
    assign memory[2255] = 16'd11269;
    assign memory[2256] = 16'd11245;
    assign memory[2257] = 16'd11221;
    assign memory[2258] = 16'd11197;
    assign memory[2259] = 16'd11174;
    assign memory[2260] = 16'd11150;
    assign memory[2261] = 16'd11126;
    assign memory[2262] = 16'd11102;
    assign memory[2263] = 16'd11078;
    assign memory[2264] = 16'd11055;
    assign memory[2265] = 16'd11031;
    assign memory[2266] = 16'd11007;
    assign memory[2267] = 16'd10983;
    assign memory[2268] = 16'd10960;
    assign memory[2269] = 16'd10936;
    assign memory[2270] = 16'd10912;
    assign memory[2271] = 16'd10889;
    assign memory[2272] = 16'd10865;
    assign memory[2273] = 16'd10841;
    assign memory[2274] = 16'd10818;
    assign memory[2275] = 16'd10794;
    assign memory[2276] = 16'd10770;
    assign memory[2277] = 16'd10747;
    assign memory[2278] = 16'd10723;
    assign memory[2279] = 16'd10700;
    assign memory[2280] = 16'd10676;
    assign memory[2281] = 16'd10652;
    assign memory[2282] = 16'd10629;
    assign memory[2283] = 16'd10605;
    assign memory[2284] = 16'd10582;
    assign memory[2285] = 16'd10558;
    assign memory[2286] = 16'd10535;
    assign memory[2287] = 16'd10511;
    assign memory[2288] = 16'd10488;
    assign memory[2289] = 16'd10465;
    assign memory[2290] = 16'd10441;
    assign memory[2291] = 16'd10418;
    assign memory[2292] = 16'd10394;
    assign memory[2293] = 16'd10371;
    assign memory[2294] = 16'd10348;
    assign memory[2295] = 16'd10324;
    assign memory[2296] = 16'd10301;
    assign memory[2297] = 16'd10278;
    assign memory[2298] = 16'd10254;
    assign memory[2299] = 16'd10231;
    assign memory[2300] = 16'd10208;
    assign memory[2301] = 16'd10184;
    assign memory[2302] = 16'd10161;
    assign memory[2303] = 16'd10138;
    assign memory[2304] = 16'd10115;
    assign memory[2305] = 16'd10091;
    assign memory[2306] = 16'd10068;
    assign memory[2307] = 16'd10045;
    assign memory[2308] = 16'd10022;
    assign memory[2309] = 16'd 9999;
    assign memory[2310] = 16'd 9976;
    assign memory[2311] = 16'd 9952;
    assign memory[2312] = 16'd 9929;
    assign memory[2313] = 16'd 9906;
    assign memory[2314] = 16'd 9883;
    assign memory[2315] = 16'd 9860;
    assign memory[2316] = 16'd 9837;
    assign memory[2317] = 16'd 9814;
    assign memory[2318] = 16'd 9791;
    assign memory[2319] = 16'd 9768;
    assign memory[2320] = 16'd 9745;
    assign memory[2321] = 16'd 9722;
    assign memory[2322] = 16'd 9699;
    assign memory[2323] = 16'd 9676;
    assign memory[2324] = 16'd 9653;
    assign memory[2325] = 16'd 9630;
    assign memory[2326] = 16'd 9607;
    assign memory[2327] = 16'd 9585;
    assign memory[2328] = 16'd 9562;
    assign memory[2329] = 16'd 9539;
    assign memory[2330] = 16'd 9516;
    assign memory[2331] = 16'd 9493;
    assign memory[2332] = 16'd 9470;
    assign memory[2333] = 16'd 9448;
    assign memory[2334] = 16'd 9425;
    assign memory[2335] = 16'd 9402;
    assign memory[2336] = 16'd 9379;
    assign memory[2337] = 16'd 9357;
    assign memory[2338] = 16'd 9334;
    assign memory[2339] = 16'd 9311;
    assign memory[2340] = 16'd 9289;
    assign memory[2341] = 16'd 9266;
    assign memory[2342] = 16'd 9243;
    assign memory[2343] = 16'd 9221;
    assign memory[2344] = 16'd 9198;
    assign memory[2345] = 16'd 9176;
    assign memory[2346] = 16'd 9153;
    assign memory[2347] = 16'd 9131;
    assign memory[2348] = 16'd 9108;
    assign memory[2349] = 16'd 9085;
    assign memory[2350] = 16'd 9063;
    assign memory[2351] = 16'd 9041;
    assign memory[2352] = 16'd 9018;
    assign memory[2353] = 16'd 8996;
    assign memory[2354] = 16'd 8973;
    assign memory[2355] = 16'd 8951;
    assign memory[2356] = 16'd 8928;
    assign memory[2357] = 16'd 8906;
    assign memory[2358] = 16'd 8884;
    assign memory[2359] = 16'd 8861;
    assign memory[2360] = 16'd 8839;
    assign memory[2361] = 16'd 8817;
    assign memory[2362] = 16'd 8794;
    assign memory[2363] = 16'd 8772;
    assign memory[2364] = 16'd 8750;
    assign memory[2365] = 16'd 8728;
    assign memory[2366] = 16'd 8706;
    assign memory[2367] = 16'd 8683;
    assign memory[2368] = 16'd 8661;
    assign memory[2369] = 16'd 8639;
    assign memory[2370] = 16'd 8617;
    assign memory[2371] = 16'd 8595;
    assign memory[2372] = 16'd 8573;
    assign memory[2373] = 16'd 8551;
    assign memory[2374] = 16'd 8528;
    assign memory[2375] = 16'd 8506;
    assign memory[2376] = 16'd 8484;
    assign memory[2377] = 16'd 8462;
    assign memory[2378] = 16'd 8440;
    assign memory[2379] = 16'd 8418;
    assign memory[2380] = 16'd 8396;
    assign memory[2381] = 16'd 8375;
    assign memory[2382] = 16'd 8353;
    assign memory[2383] = 16'd 8331;
    assign memory[2384] = 16'd 8309;
    assign memory[2385] = 16'd 8287;
    assign memory[2386] = 16'd 8265;
    assign memory[2387] = 16'd 8243;
    assign memory[2388] = 16'd 8222;
    assign memory[2389] = 16'd 8200;
    assign memory[2390] = 16'd 8178;
    assign memory[2391] = 16'd 8156;
    assign memory[2392] = 16'd 8135;
    assign memory[2393] = 16'd 8113;
    assign memory[2394] = 16'd 8091;
    assign memory[2395] = 16'd 8069;
    assign memory[2396] = 16'd 8048;
    assign memory[2397] = 16'd 8026;
    assign memory[2398] = 16'd 8005;
    assign memory[2399] = 16'd 7983;
    assign memory[2400] = 16'd 7961;
    assign memory[2401] = 16'd 7940;
    assign memory[2402] = 16'd 7918;
    assign memory[2403] = 16'd 7897;
    assign memory[2404] = 16'd 7875;
    assign memory[2405] = 16'd 7854;
    assign memory[2406] = 16'd 7832;
    assign memory[2407] = 16'd 7811;
    assign memory[2408] = 16'd 7790;
    assign memory[2409] = 16'd 7768;
    assign memory[2410] = 16'd 7747;
    assign memory[2411] = 16'd 7726;
    assign memory[2412] = 16'd 7704;
    assign memory[2413] = 16'd 7683;
    assign memory[2414] = 16'd 7662;
    assign memory[2415] = 16'd 7640;
    assign memory[2416] = 16'd 7619;
    assign memory[2417] = 16'd 7598;
    assign memory[2418] = 16'd 7577;
    assign memory[2419] = 16'd 7555;
    assign memory[2420] = 16'd 7534;
    assign memory[2421] = 16'd 7513;
    assign memory[2422] = 16'd 7492;
    assign memory[2423] = 16'd 7471;
    assign memory[2424] = 16'd 7450;
    assign memory[2425] = 16'd 7429;
    assign memory[2426] = 16'd 7408;
    assign memory[2427] = 16'd 7387;
    assign memory[2428] = 16'd 7366;
    assign memory[2429] = 16'd 7345;
    assign memory[2430] = 16'd 7324;
    assign memory[2431] = 16'd 7303;
    assign memory[2432] = 16'd 7282;
    assign memory[2433] = 16'd 7261;
    assign memory[2434] = 16'd 7240;
    assign memory[2435] = 16'd 7219;
    assign memory[2436] = 16'd 7199;
    assign memory[2437] = 16'd 7178;
    assign memory[2438] = 16'd 7157;
    assign memory[2439] = 16'd 7136;
    assign memory[2440] = 16'd 7116;
    assign memory[2441] = 16'd 7095;
    assign memory[2442] = 16'd 7074;
    assign memory[2443] = 16'd 7053;
    assign memory[2444] = 16'd 7033;
    assign memory[2445] = 16'd 7012;
    assign memory[2446] = 16'd 6992;
    assign memory[2447] = 16'd 6971;
    assign memory[2448] = 16'd 6950;
    assign memory[2449] = 16'd 6930;
    assign memory[2450] = 16'd 6909;
    assign memory[2451] = 16'd 6889;
    assign memory[2452] = 16'd 6868;
    assign memory[2453] = 16'd 6848;
    assign memory[2454] = 16'd 6828;
    assign memory[2455] = 16'd 6807;
    assign memory[2456] = 16'd 6787;
    assign memory[2457] = 16'd 6766;
    assign memory[2458] = 16'd 6746;
    assign memory[2459] = 16'd 6726;
    assign memory[2460] = 16'd 6705;
    assign memory[2461] = 16'd 6685;
    assign memory[2462] = 16'd 6665;
    assign memory[2463] = 16'd 6645;
    assign memory[2464] = 16'd 6625;
    assign memory[2465] = 16'd 6604;
    assign memory[2466] = 16'd 6584;
    assign memory[2467] = 16'd 6564;
    assign memory[2468] = 16'd 6544;
    assign memory[2469] = 16'd 6524;
    assign memory[2470] = 16'd 6504;
    assign memory[2471] = 16'd 6484;
    assign memory[2472] = 16'd 6464;
    assign memory[2473] = 16'd 6444;
    assign memory[2474] = 16'd 6424;
    assign memory[2475] = 16'd 6404;
    assign memory[2476] = 16'd 6384;
    assign memory[2477] = 16'd 6364;
    assign memory[2478] = 16'd 6344;
    assign memory[2479] = 16'd 6324;
    assign memory[2480] = 16'd 6305;
    assign memory[2481] = 16'd 6285;
    assign memory[2482] = 16'd 6265;
    assign memory[2483] = 16'd 6245;
    assign memory[2484] = 16'd 6225;
    assign memory[2485] = 16'd 6206;
    assign memory[2486] = 16'd 6186;
    assign memory[2487] = 16'd 6166;
    assign memory[2488] = 16'd 6147;
    assign memory[2489] = 16'd 6127;
    assign memory[2490] = 16'd 6108;
    assign memory[2491] = 16'd 6088;
    assign memory[2492] = 16'd 6069;
    assign memory[2493] = 16'd 6049;
    assign memory[2494] = 16'd 6030;
    assign memory[2495] = 16'd 6010;
    assign memory[2496] = 16'd 5991;
    assign memory[2497] = 16'd 5971;
    assign memory[2498] = 16'd 5952;
    assign memory[2499] = 16'd 5932;
    assign memory[2500] = 16'd 5913;
    assign memory[2501] = 16'd 5894;
    assign memory[2502] = 16'd 5874;
    assign memory[2503] = 16'd 5855;
    assign memory[2504] = 16'd 5836;
    assign memory[2505] = 16'd 5817;
    assign memory[2506] = 16'd 5798;
    assign memory[2507] = 16'd 5778;
    assign memory[2508] = 16'd 5759;
    assign memory[2509] = 16'd 5740;
    assign memory[2510] = 16'd 5721;
    assign memory[2511] = 16'd 5702;
    assign memory[2512] = 16'd 5683;
    assign memory[2513] = 16'd 5664;
    assign memory[2514] = 16'd 5645;
    assign memory[2515] = 16'd 5626;
    assign memory[2516] = 16'd 5607;
    assign memory[2517] = 16'd 5588;
    assign memory[2518] = 16'd 5569;
    assign memory[2519] = 16'd 5550;
    assign memory[2520] = 16'd 5531;
    assign memory[2521] = 16'd 5513;
    assign memory[2522] = 16'd 5494;
    assign memory[2523] = 16'd 5475;
    assign memory[2524] = 16'd 5456;
    assign memory[2525] = 16'd 5438;
    assign memory[2526] = 16'd 5419;
    assign memory[2527] = 16'd 5400;
    assign memory[2528] = 16'd 5382;
    assign memory[2529] = 16'd 5363;
    assign memory[2530] = 16'd 5344;
    assign memory[2531] = 16'd 5326;
    assign memory[2532] = 16'd 5307;
    assign memory[2533] = 16'd 5289;
    assign memory[2534] = 16'd 5270;
    assign memory[2535] = 16'd 5252;
    assign memory[2536] = 16'd 5234;
    assign memory[2537] = 16'd 5215;
    assign memory[2538] = 16'd 5197;
    assign memory[2539] = 16'd 5178;
    assign memory[2540] = 16'd 5160;
    assign memory[2541] = 16'd 5142;
    assign memory[2542] = 16'd 5124;
    assign memory[2543] = 16'd 5105;
    assign memory[2544] = 16'd 5087;
    assign memory[2545] = 16'd 5069;
    assign memory[2546] = 16'd 5051;
    assign memory[2547] = 16'd 5033;
    assign memory[2548] = 16'd 5014;
    assign memory[2549] = 16'd 4996;
    assign memory[2550] = 16'd 4978;
    assign memory[2551] = 16'd 4960;
    assign memory[2552] = 16'd 4942;
    assign memory[2553] = 16'd 4924;
    assign memory[2554] = 16'd 4906;
    assign memory[2555] = 16'd 4888;
    assign memory[2556] = 16'd 4871;
    assign memory[2557] = 16'd 4853;
    assign memory[2558] = 16'd 4835;
    assign memory[2559] = 16'd 4817;
    assign memory[2560] = 16'd 4799;
    assign memory[2561] = 16'd 4782;
    assign memory[2562] = 16'd 4764;
    assign memory[2563] = 16'd 4746;
    assign memory[2564] = 16'd 4728;
    assign memory[2565] = 16'd 4711;
    assign memory[2566] = 16'd 4693;
    assign memory[2567] = 16'd 4676;
    assign memory[2568] = 16'd 4658;
    assign memory[2569] = 16'd 4640;
    assign memory[2570] = 16'd 4623;
    assign memory[2571] = 16'd 4605;
    assign memory[2572] = 16'd 4588;
    assign memory[2573] = 16'd 4571;
    assign memory[2574] = 16'd 4553;
    assign memory[2575] = 16'd 4536;
    assign memory[2576] = 16'd 4518;
    assign memory[2577] = 16'd 4501;
    assign memory[2578] = 16'd 4484;
    assign memory[2579] = 16'd 4467;
    assign memory[2580] = 16'd 4449;
    assign memory[2581] = 16'd 4432;
    assign memory[2582] = 16'd 4415;
    assign memory[2583] = 16'd 4398;
    assign memory[2584] = 16'd 4381;
    assign memory[2585] = 16'd 4364;
    assign memory[2586] = 16'd 4347;
    assign memory[2587] = 16'd 4330;
    assign memory[2588] = 16'd 4312;
    assign memory[2589] = 16'd 4296;
    assign memory[2590] = 16'd 4279;
    assign memory[2591] = 16'd 4262;
    assign memory[2592] = 16'd 4245;
    assign memory[2593] = 16'd 4228;
    assign memory[2594] = 16'd 4211;
    assign memory[2595] = 16'd 4194;
    assign memory[2596] = 16'd 4177;
    assign memory[2597] = 16'd 4161;
    assign memory[2598] = 16'd 4144;
    assign memory[2599] = 16'd 4127;
    assign memory[2600] = 16'd 4111;
    assign memory[2601] = 16'd 4094;
    assign memory[2602] = 16'd 4077;
    assign memory[2603] = 16'd 4061;
    assign memory[2604] = 16'd 4044;
    assign memory[2605] = 16'd 4028;
    assign memory[2606] = 16'd 4011;
    assign memory[2607] = 16'd 3995;
    assign memory[2608] = 16'd 3978;
    assign memory[2609] = 16'd 3962;
    assign memory[2610] = 16'd 3946;
    assign memory[2611] = 16'd 3929;
    assign memory[2612] = 16'd 3913;
    assign memory[2613] = 16'd 3897;
    assign memory[2614] = 16'd 3880;
    assign memory[2615] = 16'd 3864;
    assign memory[2616] = 16'd 3848;
    assign memory[2617] = 16'd 3832;
    assign memory[2618] = 16'd 3816;
    assign memory[2619] = 16'd 3800;
    assign memory[2620] = 16'd 3784;
    assign memory[2621] = 16'd 3767;
    assign memory[2622] = 16'd 3751;
    assign memory[2623] = 16'd 3735;
    assign memory[2624] = 16'd 3719;
    assign memory[2625] = 16'd 3704;
    assign memory[2626] = 16'd 3688;
    assign memory[2627] = 16'd 3672;
    assign memory[2628] = 16'd 3656;
    assign memory[2629] = 16'd 3640;
    assign memory[2630] = 16'd 3624;
    assign memory[2631] = 16'd 3609;
    assign memory[2632] = 16'd 3593;
    assign memory[2633] = 16'd 3577;
    assign memory[2634] = 16'd 3562;
    assign memory[2635] = 16'd 3546;
    assign memory[2636] = 16'd 3530;
    assign memory[2637] = 16'd 3515;
    assign memory[2638] = 16'd 3499;
    assign memory[2639] = 16'd 3484;
    assign memory[2640] = 16'd 3468;
    assign memory[2641] = 16'd 3453;
    assign memory[2642] = 16'd 3437;
    assign memory[2643] = 16'd 3422;
    assign memory[2644] = 16'd 3407;
    assign memory[2645] = 16'd 3391;
    assign memory[2646] = 16'd 3376;
    assign memory[2647] = 16'd 3361;
    assign memory[2648] = 16'd 3346;
    assign memory[2649] = 16'd 3330;
    assign memory[2650] = 16'd 3315;
    assign memory[2651] = 16'd 3300;
    assign memory[2652] = 16'd 3285;
    assign memory[2653] = 16'd 3270;
    assign memory[2654] = 16'd 3255;
    assign memory[2655] = 16'd 3240;
    assign memory[2656] = 16'd 3225;
    assign memory[2657] = 16'd 3210;
    assign memory[2658] = 16'd 3195;
    assign memory[2659] = 16'd 3180;
    assign memory[2660] = 16'd 3165;
    assign memory[2661] = 16'd 3150;
    assign memory[2662] = 16'd 3135;
    assign memory[2663] = 16'd 3121;
    assign memory[2664] = 16'd 3106;
    assign memory[2665] = 16'd 3091;
    assign memory[2666] = 16'd 3077;
    assign memory[2667] = 16'd 3062;
    assign memory[2668] = 16'd 3047;
    assign memory[2669] = 16'd 3033;
    assign memory[2670] = 16'd 3018;
    assign memory[2671] = 16'd 3004;
    assign memory[2672] = 16'd 2989;
    assign memory[2673] = 16'd 2975;
    assign memory[2674] = 16'd 2960;
    assign memory[2675] = 16'd 2946;
    assign memory[2676] = 16'd 2932;
    assign memory[2677] = 16'd 2917;
    assign memory[2678] = 16'd 2903;
    assign memory[2679] = 16'd 2889;
    assign memory[2680] = 16'd 2874;
    assign memory[2681] = 16'd 2860;
    assign memory[2682] = 16'd 2846;
    assign memory[2683] = 16'd 2832;
    assign memory[2684] = 16'd 2818;
    assign memory[2685] = 16'd 2804;
    assign memory[2686] = 16'd 2790;
    assign memory[2687] = 16'd 2776;
    assign memory[2688] = 16'd 2762;
    assign memory[2689] = 16'd 2748;
    assign memory[2690] = 16'd 2734;
    assign memory[2691] = 16'd 2720;
    assign memory[2692] = 16'd 2706;
    assign memory[2693] = 16'd 2692;
    assign memory[2694] = 16'd 2679;
    assign memory[2695] = 16'd 2665;
    assign memory[2696] = 16'd 2651;
    assign memory[2697] = 16'd 2637;
    assign memory[2698] = 16'd 2624;
    assign memory[2699] = 16'd 2610;
    assign memory[2700] = 16'd 2596;
    assign memory[2701] = 16'd 2583;
    assign memory[2702] = 16'd 2569;
    assign memory[2703] = 16'd 2556;
    assign memory[2704] = 16'd 2542;
    assign memory[2705] = 16'd 2529;
    assign memory[2706] = 16'd 2516;
    assign memory[2707] = 16'd 2502;
    assign memory[2708] = 16'd 2489;
    assign memory[2709] = 16'd 2476;
    assign memory[2710] = 16'd 2462;
    assign memory[2711] = 16'd 2449;
    assign memory[2712] = 16'd 2436;
    assign memory[2713] = 16'd 2423;
    assign memory[2714] = 16'd 2410;
    assign memory[2715] = 16'd 2396;
    assign memory[2716] = 16'd 2383;
    assign memory[2717] = 16'd 2370;
    assign memory[2718] = 16'd 2357;
    assign memory[2719] = 16'd 2344;
    assign memory[2720] = 16'd 2331;
    assign memory[2721] = 16'd 2319;
    assign memory[2722] = 16'd 2306;
    assign memory[2723] = 16'd 2293;
    assign memory[2724] = 16'd 2280;
    assign memory[2725] = 16'd 2267;
    assign memory[2726] = 16'd 2255;
    assign memory[2727] = 16'd 2242;
    assign memory[2728] = 16'd 2229;
    assign memory[2729] = 16'd 2217;
    assign memory[2730] = 16'd 2204;
    assign memory[2731] = 16'd 2191;
    assign memory[2732] = 16'd 2179;
    assign memory[2733] = 16'd 2166;
    assign memory[2734] = 16'd 2154;
    assign memory[2735] = 16'd 2141;
    assign memory[2736] = 16'd 2129;
    assign memory[2737] = 16'd 2117;
    assign memory[2738] = 16'd 2104;
    assign memory[2739] = 16'd 2092;
    assign memory[2740] = 16'd 2080;
    assign memory[2741] = 16'd 2067;
    assign memory[2742] = 16'd 2055;
    assign memory[2743] = 16'd 2043;
    assign memory[2744] = 16'd 2031;
    assign memory[2745] = 16'd 2019;
    assign memory[2746] = 16'd 2007;
    assign memory[2747] = 16'd 1995;
    assign memory[2748] = 16'd 1983;
    assign memory[2749] = 16'd 1971;
    assign memory[2750] = 16'd 1959;
    assign memory[2751] = 16'd 1947;
    assign memory[2752] = 16'd 1935;
    assign memory[2753] = 16'd 1923;
    assign memory[2754] = 16'd 1911;
    assign memory[2755] = 16'd 1900;
    assign memory[2756] = 16'd 1888;
    assign memory[2757] = 16'd 1876;
    assign memory[2758] = 16'd 1865;
    assign memory[2759] = 16'd 1853;
    assign memory[2760] = 16'd 1841;
    assign memory[2761] = 16'd 1830;
    assign memory[2762] = 16'd 1818;
    assign memory[2763] = 16'd 1807;
    assign memory[2764] = 16'd 1795;
    assign memory[2765] = 16'd 1784;
    assign memory[2766] = 16'd 1773;
    assign memory[2767] = 16'd 1761;
    assign memory[2768] = 16'd 1750;
    assign memory[2769] = 16'd 1739;
    assign memory[2770] = 16'd 1727;
    assign memory[2771] = 16'd 1716;
    assign memory[2772] = 16'd 1705;
    assign memory[2773] = 16'd 1694;
    assign memory[2774] = 16'd 1683;
    assign memory[2775] = 16'd 1672;
    assign memory[2776] = 16'd 1661;
    assign memory[2777] = 16'd 1650;
    assign memory[2778] = 16'd 1639;
    assign memory[2779] = 16'd 1628;
    assign memory[2780] = 16'd 1617;
    assign memory[2781] = 16'd 1606;
    assign memory[2782] = 16'd 1595;
    assign memory[2783] = 16'd 1584;
    assign memory[2784] = 16'd 1574;
    assign memory[2785] = 16'd 1563;
    assign memory[2786] = 16'd 1552;
    assign memory[2787] = 16'd 1541;
    assign memory[2788] = 16'd 1531;
    assign memory[2789] = 16'd 1520;
    assign memory[2790] = 16'd 1510;
    assign memory[2791] = 16'd 1499;
    assign memory[2792] = 16'd 1489;
    assign memory[2793] = 16'd 1478;
    assign memory[2794] = 16'd 1468;
    assign memory[2795] = 16'd 1457;
    assign memory[2796] = 16'd 1447;
    assign memory[2797] = 16'd 1437;
    assign memory[2798] = 16'd 1427;
    assign memory[2799] = 16'd 1416;
    assign memory[2800] = 16'd 1406;
    assign memory[2801] = 16'd 1396;
    assign memory[2802] = 16'd 1386;
    assign memory[2803] = 16'd 1376;
    assign memory[2804] = 16'd 1366;
    assign memory[2805] = 16'd 1356;
    assign memory[2806] = 16'd 1346;
    assign memory[2807] = 16'd 1336;
    assign memory[2808] = 16'd 1326;
    assign memory[2809] = 16'd 1316;
    assign memory[2810] = 16'd 1306;
    assign memory[2811] = 16'd 1296;
    assign memory[2812] = 16'd 1286;
    assign memory[2813] = 16'd 1277;
    assign memory[2814] = 16'd 1267;
    assign memory[2815] = 16'd 1257;
    assign memory[2816] = 16'd 1248;
    assign memory[2817] = 16'd 1238;
    assign memory[2818] = 16'd 1228;
    assign memory[2819] = 16'd 1219;
    assign memory[2820] = 16'd 1209;
    assign memory[2821] = 16'd 1200;
    assign memory[2822] = 16'd 1191;
    assign memory[2823] = 16'd 1181;
    assign memory[2824] = 16'd 1172;
    assign memory[2825] = 16'd 1163;
    assign memory[2826] = 16'd 1153;
    assign memory[2827] = 16'd 1144;
    assign memory[2828] = 16'd 1135;
    assign memory[2829] = 16'd 1126;
    assign memory[2830] = 16'd 1117;
    assign memory[2831] = 16'd 1107;
    assign memory[2832] = 16'd 1098;
    assign memory[2833] = 16'd 1089;
    assign memory[2834] = 16'd 1080;
    assign memory[2835] = 16'd 1071;
    assign memory[2836] = 16'd 1062;
    assign memory[2837] = 16'd 1054;
    assign memory[2838] = 16'd 1045;
    assign memory[2839] = 16'd 1036;
    assign memory[2840] = 16'd 1027;
    assign memory[2841] = 16'd 1018;
    assign memory[2842] = 16'd 1010;
    assign memory[2843] = 16'd 1001;
    assign memory[2844] = 16'd  992;
    assign memory[2845] = 16'd  984;
    assign memory[2846] = 16'd  975;
    assign memory[2847] = 16'd  967;
    assign memory[2848] = 16'd  958;
    assign memory[2849] = 16'd  950;
    assign memory[2850] = 16'd  941;
    assign memory[2851] = 16'd  933;
    assign memory[2852] = 16'd  925;
    assign memory[2853] = 16'd  916;
    assign memory[2854] = 16'd  908;
    assign memory[2855] = 16'd  900;
    assign memory[2856] = 16'd  892;
    assign memory[2857] = 16'd  884;
    assign memory[2858] = 16'd  875;
    assign memory[2859] = 16'd  867;
    assign memory[2860] = 16'd  859;
    assign memory[2861] = 16'd  851;
    assign memory[2862] = 16'd  843;
    assign memory[2863] = 16'd  835;
    assign memory[2864] = 16'd  827;
    assign memory[2865] = 16'd  820;
    assign memory[2866] = 16'd  812;
    assign memory[2867] = 16'd  804;
    assign memory[2868] = 16'd  796;
    assign memory[2869] = 16'd  788;
    assign memory[2870] = 16'd  781;
    assign memory[2871] = 16'd  773;
    assign memory[2872] = 16'd  766;
    assign memory[2873] = 16'd  758;
    assign memory[2874] = 16'd  750;
    assign memory[2875] = 16'd  743;
    assign memory[2876] = 16'd  735;
    assign memory[2877] = 16'd  728;
    assign memory[2878] = 16'd  721;
    assign memory[2879] = 16'd  713;
    assign memory[2880] = 16'd  706;
    assign memory[2881] = 16'd  699;
    assign memory[2882] = 16'd  691;
    assign memory[2883] = 16'd  684;
    assign memory[2884] = 16'd  677;
    assign memory[2885] = 16'd  670;
    assign memory[2886] = 16'd  663;
    assign memory[2887] = 16'd  656;
    assign memory[2888] = 16'd  649;
    assign memory[2889] = 16'd  642;
    assign memory[2890] = 16'd  635;
    assign memory[2891] = 16'd  628;
    assign memory[2892] = 16'd  621;
    assign memory[2893] = 16'd  614;
    assign memory[2894] = 16'd  607;
    assign memory[2895] = 16'd  601;
    assign memory[2896] = 16'd  594;
    assign memory[2897] = 16'd  587;
    assign memory[2898] = 16'd  581;
    assign memory[2899] = 16'd  574;
    assign memory[2900] = 16'd  567;
    assign memory[2901] = 16'd  561;
    assign memory[2902] = 16'd  554;
    assign memory[2903] = 16'd  548;
    assign memory[2904] = 16'd  542;
    assign memory[2905] = 16'd  535;
    assign memory[2906] = 16'd  529;
    assign memory[2907] = 16'd  523;
    assign memory[2908] = 16'd  516;
    assign memory[2909] = 16'd  510;
    assign memory[2910] = 16'd  504;
    assign memory[2911] = 16'd  498;
    assign memory[2912] = 16'd  492;
    assign memory[2913] = 16'd  485;
    assign memory[2914] = 16'd  479;
    assign memory[2915] = 16'd  473;
    assign memory[2916] = 16'd  467;
    assign memory[2917] = 16'd  461;
    assign memory[2918] = 16'd  456;
    assign memory[2919] = 16'd  450;
    assign memory[2920] = 16'd  444;
    assign memory[2921] = 16'd  438;
    assign memory[2922] = 16'd  432;
    assign memory[2923] = 16'd  427;
    assign memory[2924] = 16'd  421;
    assign memory[2925] = 16'd  415;
    assign memory[2926] = 16'd  410;
    assign memory[2927] = 16'd  404;
    assign memory[2928] = 16'd  399;
    assign memory[2929] = 16'd  393;
    assign memory[2930] = 16'd  388;
    assign memory[2931] = 16'd  382;
    assign memory[2932] = 16'd  377;
    assign memory[2933] = 16'd  372;
    assign memory[2934] = 16'd  366;
    assign memory[2935] = 16'd  361;
    assign memory[2936] = 16'd  356;
    assign memory[2937] = 16'd  351;
    assign memory[2938] = 16'd  345;
    assign memory[2939] = 16'd  340;
    assign memory[2940] = 16'd  335;
    assign memory[2941] = 16'd  330;
    assign memory[2942] = 16'd  325;
    assign memory[2943] = 16'd  320;
    assign memory[2944] = 16'd  315;
    assign memory[2945] = 16'd  310;
    assign memory[2946] = 16'd  306;
    assign memory[2947] = 16'd  301;
    assign memory[2948] = 16'd  296;
    assign memory[2949] = 16'd  291;
    assign memory[2950] = 16'd  287;
    assign memory[2951] = 16'd  282;
    assign memory[2952] = 16'd  277;
    assign memory[2953] = 16'd  273;
    assign memory[2954] = 16'd  268;
    assign memory[2955] = 16'd  264;
    assign memory[2956] = 16'd  259;
    assign memory[2957] = 16'd  255;
    assign memory[2958] = 16'd  250;
    assign memory[2959] = 16'd  246;
    assign memory[2960] = 16'd  242;
    assign memory[2961] = 16'd  237;
    assign memory[2962] = 16'd  233;
    assign memory[2963] = 16'd  229;
    assign memory[2964] = 16'd  225;
    assign memory[2965] = 16'd  221;
    assign memory[2966] = 16'd  217;
    assign memory[2967] = 16'd  213;
    assign memory[2968] = 16'd  209;
    assign memory[2969] = 16'd  205;
    assign memory[2970] = 16'd  201;
    assign memory[2971] = 16'd  197;
    assign memory[2972] = 16'd  193;
    assign memory[2973] = 16'd  189;
    assign memory[2974] = 16'd  185;
    assign memory[2975] = 16'd  182;
    assign memory[2976] = 16'd  178;
    assign memory[2977] = 16'd  174;
    assign memory[2978] = 16'd  171;
    assign memory[2979] = 16'd  167;
    assign memory[2980] = 16'd  163;
    assign memory[2981] = 16'd  160;
    assign memory[2982] = 16'd  156;
    assign memory[2983] = 16'd  153;
    assign memory[2984] = 16'd  150;
    assign memory[2985] = 16'd  146;
    assign memory[2986] = 16'd  143;
    assign memory[2987] = 16'd  140;
    assign memory[2988] = 16'd  136;
    assign memory[2989] = 16'd  133;
    assign memory[2990] = 16'd  130;
    assign memory[2991] = 16'd  127;
    assign memory[2992] = 16'd  124;
    assign memory[2993] = 16'd  121;
    assign memory[2994] = 16'd  118;
    assign memory[2995] = 16'd  115;
    assign memory[2996] = 16'd  112;
    assign memory[2997] = 16'd  109;
    assign memory[2998] = 16'd  106;
    assign memory[2999] = 16'd  103;
    assign memory[3000] = 16'd  100;
    assign memory[3001] = 16'd   98;
    assign memory[3002] = 16'd   95;
    assign memory[3003] = 16'd   92;
    assign memory[3004] = 16'd   90;
    assign memory[3005] = 16'd   87;
    assign memory[3006] = 16'd   84;
    assign memory[3007] = 16'd   82;
    assign memory[3008] = 16'd   79;
    assign memory[3009] = 16'd   77;
    assign memory[3010] = 16'd   75;
    assign memory[3011] = 16'd   72;
    assign memory[3012] = 16'd   70;
    assign memory[3013] = 16'd   68;
    assign memory[3014] = 16'd   65;
    assign memory[3015] = 16'd   63;
    assign memory[3016] = 16'd   61;
    assign memory[3017] = 16'd   59;
    assign memory[3018] = 16'd   57;
    assign memory[3019] = 16'd   55;
    assign memory[3020] = 16'd   53;
    assign memory[3021] = 16'd   51;
    assign memory[3022] = 16'd   49;
    assign memory[3023] = 16'd   47;
    assign memory[3024] = 16'd   45;
    assign memory[3025] = 16'd   43;
    assign memory[3026] = 16'd   41;
    assign memory[3027] = 16'd   40;
    assign memory[3028] = 16'd   38;
    assign memory[3029] = 16'd   36;
    assign memory[3030] = 16'd   34;
    assign memory[3031] = 16'd   33;
    assign memory[3032] = 16'd   31;
    assign memory[3033] = 16'd   30;
    assign memory[3034] = 16'd   28;
    assign memory[3035] = 16'd   27;
    assign memory[3036] = 16'd   25;
    assign memory[3037] = 16'd   24;
    assign memory[3038] = 16'd   23;
    assign memory[3039] = 16'd   21;
    assign memory[3040] = 16'd   20;
    assign memory[3041] = 16'd   19;
    assign memory[3042] = 16'd   18;
    assign memory[3043] = 16'd   17;
    assign memory[3044] = 16'd   16;
    assign memory[3045] = 16'd   15;
    assign memory[3046] = 16'd   14;
    assign memory[3047] = 16'd   13;
    assign memory[3048] = 16'd   12;
    assign memory[3049] = 16'd   11;
    assign memory[3050] = 16'd   10;
    assign memory[3051] = 16'd    9;
    assign memory[3052] = 16'd    8;
    assign memory[3053] = 16'd    7;
    assign memory[3054] = 16'd    7;
    assign memory[3055] = 16'd    6;
    assign memory[3056] = 16'd    5;
    assign memory[3057] = 16'd    5;
    assign memory[3058] = 16'd    4;
    assign memory[3059] = 16'd    4;
    assign memory[3060] = 16'd    3;
    assign memory[3061] = 16'd    3;
    assign memory[3062] = 16'd    2;
    assign memory[3063] = 16'd    2;
    assign memory[3064] = 16'd    2;
    assign memory[3065] = 16'd    1;
    assign memory[3066] = 16'd    1;
    assign memory[3067] = 16'd    1;
    assign memory[3068] = 16'd    1;
    assign memory[3069] = 16'd    1;
    assign memory[3070] = 16'd    1;
    assign memory[3071] = 16'd    1;
    assign memory[3072] = 16'd    0;
    assign memory[3073] = 16'd    1;
    assign memory[3074] = 16'd    1;
    assign memory[3075] = 16'd    1;
    assign memory[3076] = 16'd    1;
    assign memory[3077] = 16'd    1;
    assign memory[3078] = 16'd    1;
    assign memory[3079] = 16'd    1;
    assign memory[3080] = 16'd    2;
    assign memory[3081] = 16'd    2;
    assign memory[3082] = 16'd    2;
    assign memory[3083] = 16'd    3;
    assign memory[3084] = 16'd    3;
    assign memory[3085] = 16'd    4;
    assign memory[3086] = 16'd    4;
    assign memory[3087] = 16'd    5;
    assign memory[3088] = 16'd    5;
    assign memory[3089] = 16'd    6;
    assign memory[3090] = 16'd    7;
    assign memory[3091] = 16'd    7;
    assign memory[3092] = 16'd    8;
    assign memory[3093] = 16'd    9;
    assign memory[3094] = 16'd   10;
    assign memory[3095] = 16'd   11;
    assign memory[3096] = 16'd   12;
    assign memory[3097] = 16'd   13;
    assign memory[3098] = 16'd   14;
    assign memory[3099] = 16'd   15;
    assign memory[3100] = 16'd   16;
    assign memory[3101] = 16'd   17;
    assign memory[3102] = 16'd   18;
    assign memory[3103] = 16'd   19;
    assign memory[3104] = 16'd   20;
    assign memory[3105] = 16'd   21;
    assign memory[3106] = 16'd   23;
    assign memory[3107] = 16'd   24;
    assign memory[3108] = 16'd   25;
    assign memory[3109] = 16'd   27;
    assign memory[3110] = 16'd   28;
    assign memory[3111] = 16'd   30;
    assign memory[3112] = 16'd   31;
    assign memory[3113] = 16'd   33;
    assign memory[3114] = 16'd   34;
    assign memory[3115] = 16'd   36;
    assign memory[3116] = 16'd   38;
    assign memory[3117] = 16'd   40;
    assign memory[3118] = 16'd   41;
    assign memory[3119] = 16'd   43;
    assign memory[3120] = 16'd   45;
    assign memory[3121] = 16'd   47;
    assign memory[3122] = 16'd   49;
    assign memory[3123] = 16'd   51;
    assign memory[3124] = 16'd   53;
    assign memory[3125] = 16'd   55;
    assign memory[3126] = 16'd   57;
    assign memory[3127] = 16'd   59;
    assign memory[3128] = 16'd   61;
    assign memory[3129] = 16'd   63;
    assign memory[3130] = 16'd   65;
    assign memory[3131] = 16'd   68;
    assign memory[3132] = 16'd   70;
    assign memory[3133] = 16'd   72;
    assign memory[3134] = 16'd   75;
    assign memory[3135] = 16'd   77;
    assign memory[3136] = 16'd   79;
    assign memory[3137] = 16'd   82;
    assign memory[3138] = 16'd   84;
    assign memory[3139] = 16'd   87;
    assign memory[3140] = 16'd   90;
    assign memory[3141] = 16'd   92;
    assign memory[3142] = 16'd   95;
    assign memory[3143] = 16'd   98;
    assign memory[3144] = 16'd  100;
    assign memory[3145] = 16'd  103;
    assign memory[3146] = 16'd  106;
    assign memory[3147] = 16'd  109;
    assign memory[3148] = 16'd  112;
    assign memory[3149] = 16'd  115;
    assign memory[3150] = 16'd  118;
    assign memory[3151] = 16'd  121;
    assign memory[3152] = 16'd  124;
    assign memory[3153] = 16'd  127;
    assign memory[3154] = 16'd  130;
    assign memory[3155] = 16'd  133;
    assign memory[3156] = 16'd  136;
    assign memory[3157] = 16'd  140;
    assign memory[3158] = 16'd  143;
    assign memory[3159] = 16'd  146;
    assign memory[3160] = 16'd  150;
    assign memory[3161] = 16'd  153;
    assign memory[3162] = 16'd  156;
    assign memory[3163] = 16'd  160;
    assign memory[3164] = 16'd  163;
    assign memory[3165] = 16'd  167;
    assign memory[3166] = 16'd  171;
    assign memory[3167] = 16'd  174;
    assign memory[3168] = 16'd  178;
    assign memory[3169] = 16'd  182;
    assign memory[3170] = 16'd  185;
    assign memory[3171] = 16'd  189;
    assign memory[3172] = 16'd  193;
    assign memory[3173] = 16'd  197;
    assign memory[3174] = 16'd  201;
    assign memory[3175] = 16'd  205;
    assign memory[3176] = 16'd  209;
    assign memory[3177] = 16'd  213;
    assign memory[3178] = 16'd  217;
    assign memory[3179] = 16'd  221;
    assign memory[3180] = 16'd  225;
    assign memory[3181] = 16'd  229;
    assign memory[3182] = 16'd  233;
    assign memory[3183] = 16'd  237;
    assign memory[3184] = 16'd  242;
    assign memory[3185] = 16'd  246;
    assign memory[3186] = 16'd  250;
    assign memory[3187] = 16'd  255;
    assign memory[3188] = 16'd  259;
    assign memory[3189] = 16'd  264;
    assign memory[3190] = 16'd  268;
    assign memory[3191] = 16'd  273;
    assign memory[3192] = 16'd  277;
    assign memory[3193] = 16'd  282;
    assign memory[3194] = 16'd  287;
    assign memory[3195] = 16'd  291;
    assign memory[3196] = 16'd  296;
    assign memory[3197] = 16'd  301;
    assign memory[3198] = 16'd  306;
    assign memory[3199] = 16'd  310;
    assign memory[3200] = 16'd  315;
    assign memory[3201] = 16'd  320;
    assign memory[3202] = 16'd  325;
    assign memory[3203] = 16'd  330;
    assign memory[3204] = 16'd  335;
    assign memory[3205] = 16'd  340;
    assign memory[3206] = 16'd  345;
    assign memory[3207] = 16'd  351;
    assign memory[3208] = 16'd  356;
    assign memory[3209] = 16'd  361;
    assign memory[3210] = 16'd  366;
    assign memory[3211] = 16'd  372;
    assign memory[3212] = 16'd  377;
    assign memory[3213] = 16'd  382;
    assign memory[3214] = 16'd  388;
    assign memory[3215] = 16'd  393;
    assign memory[3216] = 16'd  399;
    assign memory[3217] = 16'd  404;
    assign memory[3218] = 16'd  410;
    assign memory[3219] = 16'd  415;
    assign memory[3220] = 16'd  421;
    assign memory[3221] = 16'd  427;
    assign memory[3222] = 16'd  432;
    assign memory[3223] = 16'd  438;
    assign memory[3224] = 16'd  444;
    assign memory[3225] = 16'd  450;
    assign memory[3226] = 16'd  456;
    assign memory[3227] = 16'd  461;
    assign memory[3228] = 16'd  467;
    assign memory[3229] = 16'd  473;
    assign memory[3230] = 16'd  479;
    assign memory[3231] = 16'd  485;
    assign memory[3232] = 16'd  492;
    assign memory[3233] = 16'd  498;
    assign memory[3234] = 16'd  504;
    assign memory[3235] = 16'd  510;
    assign memory[3236] = 16'd  516;
    assign memory[3237] = 16'd  523;
    assign memory[3238] = 16'd  529;
    assign memory[3239] = 16'd  535;
    assign memory[3240] = 16'd  542;
    assign memory[3241] = 16'd  548;
    assign memory[3242] = 16'd  554;
    assign memory[3243] = 16'd  561;
    assign memory[3244] = 16'd  567;
    assign memory[3245] = 16'd  574;
    assign memory[3246] = 16'd  581;
    assign memory[3247] = 16'd  587;
    assign memory[3248] = 16'd  594;
    assign memory[3249] = 16'd  601;
    assign memory[3250] = 16'd  607;
    assign memory[3251] = 16'd  614;
    assign memory[3252] = 16'd  621;
    assign memory[3253] = 16'd  628;
    assign memory[3254] = 16'd  635;
    assign memory[3255] = 16'd  642;
    assign memory[3256] = 16'd  649;
    assign memory[3257] = 16'd  656;
    assign memory[3258] = 16'd  663;
    assign memory[3259] = 16'd  670;
    assign memory[3260] = 16'd  677;
    assign memory[3261] = 16'd  684;
    assign memory[3262] = 16'd  691;
    assign memory[3263] = 16'd  699;
    assign memory[3264] = 16'd  706;
    assign memory[3265] = 16'd  713;
    assign memory[3266] = 16'd  721;
    assign memory[3267] = 16'd  728;
    assign memory[3268] = 16'd  735;
    assign memory[3269] = 16'd  743;
    assign memory[3270] = 16'd  750;
    assign memory[3271] = 16'd  758;
    assign memory[3272] = 16'd  766;
    assign memory[3273] = 16'd  773;
    assign memory[3274] = 16'd  781;
    assign memory[3275] = 16'd  788;
    assign memory[3276] = 16'd  796;
    assign memory[3277] = 16'd  804;
    assign memory[3278] = 16'd  812;
    assign memory[3279] = 16'd  820;
    assign memory[3280] = 16'd  827;
    assign memory[3281] = 16'd  835;
    assign memory[3282] = 16'd  843;
    assign memory[3283] = 16'd  851;
    assign memory[3284] = 16'd  859;
    assign memory[3285] = 16'd  867;
    assign memory[3286] = 16'd  875;
    assign memory[3287] = 16'd  884;
    assign memory[3288] = 16'd  892;
    assign memory[3289] = 16'd  900;
    assign memory[3290] = 16'd  908;
    assign memory[3291] = 16'd  916;
    assign memory[3292] = 16'd  925;
    assign memory[3293] = 16'd  933;
    assign memory[3294] = 16'd  941;
    assign memory[3295] = 16'd  950;
    assign memory[3296] = 16'd  958;
    assign memory[3297] = 16'd  967;
    assign memory[3298] = 16'd  975;
    assign memory[3299] = 16'd  984;
    assign memory[3300] = 16'd  992;
    assign memory[3301] = 16'd 1001;
    assign memory[3302] = 16'd 1010;
    assign memory[3303] = 16'd 1018;
    assign memory[3304] = 16'd 1027;
    assign memory[3305] = 16'd 1036;
    assign memory[3306] = 16'd 1045;
    assign memory[3307] = 16'd 1054;
    assign memory[3308] = 16'd 1062;
    assign memory[3309] = 16'd 1071;
    assign memory[3310] = 16'd 1080;
    assign memory[3311] = 16'd 1089;
    assign memory[3312] = 16'd 1098;
    assign memory[3313] = 16'd 1107;
    assign memory[3314] = 16'd 1117;
    assign memory[3315] = 16'd 1126;
    assign memory[3316] = 16'd 1135;
    assign memory[3317] = 16'd 1144;
    assign memory[3318] = 16'd 1153;
    assign memory[3319] = 16'd 1163;
    assign memory[3320] = 16'd 1172;
    assign memory[3321] = 16'd 1181;
    assign memory[3322] = 16'd 1191;
    assign memory[3323] = 16'd 1200;
    assign memory[3324] = 16'd 1209;
    assign memory[3325] = 16'd 1219;
    assign memory[3326] = 16'd 1228;
    assign memory[3327] = 16'd 1238;
    assign memory[3328] = 16'd 1248;
    assign memory[3329] = 16'd 1257;
    assign memory[3330] = 16'd 1267;
    assign memory[3331] = 16'd 1277;
    assign memory[3332] = 16'd 1286;
    assign memory[3333] = 16'd 1296;
    assign memory[3334] = 16'd 1306;
    assign memory[3335] = 16'd 1316;
    assign memory[3336] = 16'd 1326;
    assign memory[3337] = 16'd 1336;
    assign memory[3338] = 16'd 1346;
    assign memory[3339] = 16'd 1356;
    assign memory[3340] = 16'd 1366;
    assign memory[3341] = 16'd 1376;
    assign memory[3342] = 16'd 1386;
    assign memory[3343] = 16'd 1396;
    assign memory[3344] = 16'd 1406;
    assign memory[3345] = 16'd 1416;
    assign memory[3346] = 16'd 1427;
    assign memory[3347] = 16'd 1437;
    assign memory[3348] = 16'd 1447;
    assign memory[3349] = 16'd 1457;
    assign memory[3350] = 16'd 1468;
    assign memory[3351] = 16'd 1478;
    assign memory[3352] = 16'd 1489;
    assign memory[3353] = 16'd 1499;
    assign memory[3354] = 16'd 1510;
    assign memory[3355] = 16'd 1520;
    assign memory[3356] = 16'd 1531;
    assign memory[3357] = 16'd 1541;
    assign memory[3358] = 16'd 1552;
    assign memory[3359] = 16'd 1563;
    assign memory[3360] = 16'd 1574;
    assign memory[3361] = 16'd 1584;
    assign memory[3362] = 16'd 1595;
    assign memory[3363] = 16'd 1606;
    assign memory[3364] = 16'd 1617;
    assign memory[3365] = 16'd 1628;
    assign memory[3366] = 16'd 1639;
    assign memory[3367] = 16'd 1650;
    assign memory[3368] = 16'd 1661;
    assign memory[3369] = 16'd 1672;
    assign memory[3370] = 16'd 1683;
    assign memory[3371] = 16'd 1694;
    assign memory[3372] = 16'd 1705;
    assign memory[3373] = 16'd 1716;
    assign memory[3374] = 16'd 1727;
    assign memory[3375] = 16'd 1739;
    assign memory[3376] = 16'd 1750;
    assign memory[3377] = 16'd 1761;
    assign memory[3378] = 16'd 1773;
    assign memory[3379] = 16'd 1784;
    assign memory[3380] = 16'd 1795;
    assign memory[3381] = 16'd 1807;
    assign memory[3382] = 16'd 1818;
    assign memory[3383] = 16'd 1830;
    assign memory[3384] = 16'd 1841;
    assign memory[3385] = 16'd 1853;
    assign memory[3386] = 16'd 1865;
    assign memory[3387] = 16'd 1876;
    assign memory[3388] = 16'd 1888;
    assign memory[3389] = 16'd 1900;
    assign memory[3390] = 16'd 1911;
    assign memory[3391] = 16'd 1923;
    assign memory[3392] = 16'd 1935;
    assign memory[3393] = 16'd 1947;
    assign memory[3394] = 16'd 1959;
    assign memory[3395] = 16'd 1971;
    assign memory[3396] = 16'd 1983;
    assign memory[3397] = 16'd 1995;
    assign memory[3398] = 16'd 2007;
    assign memory[3399] = 16'd 2019;
    assign memory[3400] = 16'd 2031;
    assign memory[3401] = 16'd 2043;
    assign memory[3402] = 16'd 2055;
    assign memory[3403] = 16'd 2067;
    assign memory[3404] = 16'd 2080;
    assign memory[3405] = 16'd 2092;
    assign memory[3406] = 16'd 2104;
    assign memory[3407] = 16'd 2117;
    assign memory[3408] = 16'd 2129;
    assign memory[3409] = 16'd 2141;
    assign memory[3410] = 16'd 2154;
    assign memory[3411] = 16'd 2166;
    assign memory[3412] = 16'd 2179;
    assign memory[3413] = 16'd 2191;
    assign memory[3414] = 16'd 2204;
    assign memory[3415] = 16'd 2217;
    assign memory[3416] = 16'd 2229;
    assign memory[3417] = 16'd 2242;
    assign memory[3418] = 16'd 2255;
    assign memory[3419] = 16'd 2267;
    assign memory[3420] = 16'd 2280;
    assign memory[3421] = 16'd 2293;
    assign memory[3422] = 16'd 2306;
    assign memory[3423] = 16'd 2319;
    assign memory[3424] = 16'd 2331;
    assign memory[3425] = 16'd 2344;
    assign memory[3426] = 16'd 2357;
    assign memory[3427] = 16'd 2370;
    assign memory[3428] = 16'd 2383;
    assign memory[3429] = 16'd 2396;
    assign memory[3430] = 16'd 2410;
    assign memory[3431] = 16'd 2423;
    assign memory[3432] = 16'd 2436;
    assign memory[3433] = 16'd 2449;
    assign memory[3434] = 16'd 2462;
    assign memory[3435] = 16'd 2476;
    assign memory[3436] = 16'd 2489;
    assign memory[3437] = 16'd 2502;
    assign memory[3438] = 16'd 2516;
    assign memory[3439] = 16'd 2529;
    assign memory[3440] = 16'd 2542;
    assign memory[3441] = 16'd 2556;
    assign memory[3442] = 16'd 2569;
    assign memory[3443] = 16'd 2583;
    assign memory[3444] = 16'd 2596;
    assign memory[3445] = 16'd 2610;
    assign memory[3446] = 16'd 2624;
    assign memory[3447] = 16'd 2637;
    assign memory[3448] = 16'd 2651;
    assign memory[3449] = 16'd 2665;
    assign memory[3450] = 16'd 2679;
    assign memory[3451] = 16'd 2692;
    assign memory[3452] = 16'd 2706;
    assign memory[3453] = 16'd 2720;
    assign memory[3454] = 16'd 2734;
    assign memory[3455] = 16'd 2748;
    assign memory[3456] = 16'd 2762;
    assign memory[3457] = 16'd 2776;
    assign memory[3458] = 16'd 2790;
    assign memory[3459] = 16'd 2804;
    assign memory[3460] = 16'd 2818;
    assign memory[3461] = 16'd 2832;
    assign memory[3462] = 16'd 2846;
    assign memory[3463] = 16'd 2860;
    assign memory[3464] = 16'd 2874;
    assign memory[3465] = 16'd 2889;
    assign memory[3466] = 16'd 2903;
    assign memory[3467] = 16'd 2917;
    assign memory[3468] = 16'd 2932;
    assign memory[3469] = 16'd 2946;
    assign memory[3470] = 16'd 2960;
    assign memory[3471] = 16'd 2975;
    assign memory[3472] = 16'd 2989;
    assign memory[3473] = 16'd 3004;
    assign memory[3474] = 16'd 3018;
    assign memory[3475] = 16'd 3033;
    assign memory[3476] = 16'd 3047;
    assign memory[3477] = 16'd 3062;
    assign memory[3478] = 16'd 3077;
    assign memory[3479] = 16'd 3091;
    assign memory[3480] = 16'd 3106;
    assign memory[3481] = 16'd 3121;
    assign memory[3482] = 16'd 3135;
    assign memory[3483] = 16'd 3150;
    assign memory[3484] = 16'd 3165;
    assign memory[3485] = 16'd 3180;
    assign memory[3486] = 16'd 3195;
    assign memory[3487] = 16'd 3210;
    assign memory[3488] = 16'd 3225;
    assign memory[3489] = 16'd 3240;
    assign memory[3490] = 16'd 3255;
    assign memory[3491] = 16'd 3270;
    assign memory[3492] = 16'd 3285;
    assign memory[3493] = 16'd 3300;
    assign memory[3494] = 16'd 3315;
    assign memory[3495] = 16'd 3330;
    assign memory[3496] = 16'd 3346;
    assign memory[3497] = 16'd 3361;
    assign memory[3498] = 16'd 3376;
    assign memory[3499] = 16'd 3391;
    assign memory[3500] = 16'd 3407;
    assign memory[3501] = 16'd 3422;
    assign memory[3502] = 16'd 3437;
    assign memory[3503] = 16'd 3453;
    assign memory[3504] = 16'd 3468;
    assign memory[3505] = 16'd 3484;
    assign memory[3506] = 16'd 3499;
    assign memory[3507] = 16'd 3515;
    assign memory[3508] = 16'd 3530;
    assign memory[3509] = 16'd 3546;
    assign memory[3510] = 16'd 3562;
    assign memory[3511] = 16'd 3577;
    assign memory[3512] = 16'd 3593;
    assign memory[3513] = 16'd 3609;
    assign memory[3514] = 16'd 3624;
    assign memory[3515] = 16'd 3640;
    assign memory[3516] = 16'd 3656;
    assign memory[3517] = 16'd 3672;
    assign memory[3518] = 16'd 3688;
    assign memory[3519] = 16'd 3704;
    assign memory[3520] = 16'd 3719;
    assign memory[3521] = 16'd 3735;
    assign memory[3522] = 16'd 3751;
    assign memory[3523] = 16'd 3767;
    assign memory[3524] = 16'd 3784;
    assign memory[3525] = 16'd 3800;
    assign memory[3526] = 16'd 3816;
    assign memory[3527] = 16'd 3832;
    assign memory[3528] = 16'd 3848;
    assign memory[3529] = 16'd 3864;
    assign memory[3530] = 16'd 3880;
    assign memory[3531] = 16'd 3897;
    assign memory[3532] = 16'd 3913;
    assign memory[3533] = 16'd 3929;
    assign memory[3534] = 16'd 3946;
    assign memory[3535] = 16'd 3962;
    assign memory[3536] = 16'd 3978;
    assign memory[3537] = 16'd 3995;
    assign memory[3538] = 16'd 4011;
    assign memory[3539] = 16'd 4028;
    assign memory[3540] = 16'd 4044;
    assign memory[3541] = 16'd 4061;
    assign memory[3542] = 16'd 4077;
    assign memory[3543] = 16'd 4094;
    assign memory[3544] = 16'd 4111;
    assign memory[3545] = 16'd 4127;
    assign memory[3546] = 16'd 4144;
    assign memory[3547] = 16'd 4161;
    assign memory[3548] = 16'd 4177;
    assign memory[3549] = 16'd 4194;
    assign memory[3550] = 16'd 4211;
    assign memory[3551] = 16'd 4228;
    assign memory[3552] = 16'd 4245;
    assign memory[3553] = 16'd 4262;
    assign memory[3554] = 16'd 4279;
    assign memory[3555] = 16'd 4296;
    assign memory[3556] = 16'd 4312;
    assign memory[3557] = 16'd 4330;
    assign memory[3558] = 16'd 4347;
    assign memory[3559] = 16'd 4364;
    assign memory[3560] = 16'd 4381;
    assign memory[3561] = 16'd 4398;
    assign memory[3562] = 16'd 4415;
    assign memory[3563] = 16'd 4432;
    assign memory[3564] = 16'd 4449;
    assign memory[3565] = 16'd 4467;
    assign memory[3566] = 16'd 4484;
    assign memory[3567] = 16'd 4501;
    assign memory[3568] = 16'd 4518;
    assign memory[3569] = 16'd 4536;
    assign memory[3570] = 16'd 4553;
    assign memory[3571] = 16'd 4571;
    assign memory[3572] = 16'd 4588;
    assign memory[3573] = 16'd 4605;
    assign memory[3574] = 16'd 4623;
    assign memory[3575] = 16'd 4640;
    assign memory[3576] = 16'd 4658;
    assign memory[3577] = 16'd 4676;
    assign memory[3578] = 16'd 4693;
    assign memory[3579] = 16'd 4711;
    assign memory[3580] = 16'd 4728;
    assign memory[3581] = 16'd 4746;
    assign memory[3582] = 16'd 4764;
    assign memory[3583] = 16'd 4782;
    assign memory[3584] = 16'd 4799;
    assign memory[3585] = 16'd 4817;
    assign memory[3586] = 16'd 4835;
    assign memory[3587] = 16'd 4853;
    assign memory[3588] = 16'd 4871;
    assign memory[3589] = 16'd 4888;
    assign memory[3590] = 16'd 4906;
    assign memory[3591] = 16'd 4924;
    assign memory[3592] = 16'd 4942;
    assign memory[3593] = 16'd 4960;
    assign memory[3594] = 16'd 4978;
    assign memory[3595] = 16'd 4996;
    assign memory[3596] = 16'd 5014;
    assign memory[3597] = 16'd 5033;
    assign memory[3598] = 16'd 5051;
    assign memory[3599] = 16'd 5069;
    assign memory[3600] = 16'd 5087;
    assign memory[3601] = 16'd 5105;
    assign memory[3602] = 16'd 5124;
    assign memory[3603] = 16'd 5142;
    assign memory[3604] = 16'd 5160;
    assign memory[3605] = 16'd 5178;
    assign memory[3606] = 16'd 5197;
    assign memory[3607] = 16'd 5215;
    assign memory[3608] = 16'd 5234;
    assign memory[3609] = 16'd 5252;
    assign memory[3610] = 16'd 5270;
    assign memory[3611] = 16'd 5289;
    assign memory[3612] = 16'd 5307;
    assign memory[3613] = 16'd 5326;
    assign memory[3614] = 16'd 5344;
    assign memory[3615] = 16'd 5363;
    assign memory[3616] = 16'd 5382;
    assign memory[3617] = 16'd 5400;
    assign memory[3618] = 16'd 5419;
    assign memory[3619] = 16'd 5438;
    assign memory[3620] = 16'd 5456;
    assign memory[3621] = 16'd 5475;
    assign memory[3622] = 16'd 5494;
    assign memory[3623] = 16'd 5513;
    assign memory[3624] = 16'd 5531;
    assign memory[3625] = 16'd 5550;
    assign memory[3626] = 16'd 5569;
    assign memory[3627] = 16'd 5588;
    assign memory[3628] = 16'd 5607;
    assign memory[3629] = 16'd 5626;
    assign memory[3630] = 16'd 5645;
    assign memory[3631] = 16'd 5664;
    assign memory[3632] = 16'd 5683;
    assign memory[3633] = 16'd 5702;
    assign memory[3634] = 16'd 5721;
    assign memory[3635] = 16'd 5740;
    assign memory[3636] = 16'd 5759;
    assign memory[3637] = 16'd 5778;
    assign memory[3638] = 16'd 5798;
    assign memory[3639] = 16'd 5817;
    assign memory[3640] = 16'd 5836;
    assign memory[3641] = 16'd 5855;
    assign memory[3642] = 16'd 5874;
    assign memory[3643] = 16'd 5894;
    assign memory[3644] = 16'd 5913;
    assign memory[3645] = 16'd 5932;
    assign memory[3646] = 16'd 5952;
    assign memory[3647] = 16'd 5971;
    assign memory[3648] = 16'd 5991;
    assign memory[3649] = 16'd 6010;
    assign memory[3650] = 16'd 6030;
    assign memory[3651] = 16'd 6049;
    assign memory[3652] = 16'd 6069;
    assign memory[3653] = 16'd 6088;
    assign memory[3654] = 16'd 6108;
    assign memory[3655] = 16'd 6127;
    assign memory[3656] = 16'd 6147;
    assign memory[3657] = 16'd 6166;
    assign memory[3658] = 16'd 6186;
    assign memory[3659] = 16'd 6206;
    assign memory[3660] = 16'd 6225;
    assign memory[3661] = 16'd 6245;
    assign memory[3662] = 16'd 6265;
    assign memory[3663] = 16'd 6285;
    assign memory[3664] = 16'd 6305;
    assign memory[3665] = 16'd 6324;
    assign memory[3666] = 16'd 6344;
    assign memory[3667] = 16'd 6364;
    assign memory[3668] = 16'd 6384;
    assign memory[3669] = 16'd 6404;
    assign memory[3670] = 16'd 6424;
    assign memory[3671] = 16'd 6444;
    assign memory[3672] = 16'd 6464;
    assign memory[3673] = 16'd 6484;
    assign memory[3674] = 16'd 6504;
    assign memory[3675] = 16'd 6524;
    assign memory[3676] = 16'd 6544;
    assign memory[3677] = 16'd 6564;
    assign memory[3678] = 16'd 6584;
    assign memory[3679] = 16'd 6604;
    assign memory[3680] = 16'd 6625;
    assign memory[3681] = 16'd 6645;
    assign memory[3682] = 16'd 6665;
    assign memory[3683] = 16'd 6685;
    assign memory[3684] = 16'd 6705;
    assign memory[3685] = 16'd 6726;
    assign memory[3686] = 16'd 6746;
    assign memory[3687] = 16'd 6766;
    assign memory[3688] = 16'd 6787;
    assign memory[3689] = 16'd 6807;
    assign memory[3690] = 16'd 6828;
    assign memory[3691] = 16'd 6848;
    assign memory[3692] = 16'd 6868;
    assign memory[3693] = 16'd 6889;
    assign memory[3694] = 16'd 6909;
    assign memory[3695] = 16'd 6930;
    assign memory[3696] = 16'd 6950;
    assign memory[3697] = 16'd 6971;
    assign memory[3698] = 16'd 6992;
    assign memory[3699] = 16'd 7012;
    assign memory[3700] = 16'd 7033;
    assign memory[3701] = 16'd 7053;
    assign memory[3702] = 16'd 7074;
    assign memory[3703] = 16'd 7095;
    assign memory[3704] = 16'd 7116;
    assign memory[3705] = 16'd 7136;
    assign memory[3706] = 16'd 7157;
    assign memory[3707] = 16'd 7178;
    assign memory[3708] = 16'd 7199;
    assign memory[3709] = 16'd 7219;
    assign memory[3710] = 16'd 7240;
    assign memory[3711] = 16'd 7261;
    assign memory[3712] = 16'd 7282;
    assign memory[3713] = 16'd 7303;
    assign memory[3714] = 16'd 7324;
    assign memory[3715] = 16'd 7345;
    assign memory[3716] = 16'd 7366;
    assign memory[3717] = 16'd 7387;
    assign memory[3718] = 16'd 7408;
    assign memory[3719] = 16'd 7429;
    assign memory[3720] = 16'd 7450;
    assign memory[3721] = 16'd 7471;
    assign memory[3722] = 16'd 7492;
    assign memory[3723] = 16'd 7513;
    assign memory[3724] = 16'd 7534;
    assign memory[3725] = 16'd 7555;
    assign memory[3726] = 16'd 7577;
    assign memory[3727] = 16'd 7598;
    assign memory[3728] = 16'd 7619;
    assign memory[3729] = 16'd 7640;
    assign memory[3730] = 16'd 7662;
    assign memory[3731] = 16'd 7683;
    assign memory[3732] = 16'd 7704;
    assign memory[3733] = 16'd 7726;
    assign memory[3734] = 16'd 7747;
    assign memory[3735] = 16'd 7768;
    assign memory[3736] = 16'd 7790;
    assign memory[3737] = 16'd 7811;
    assign memory[3738] = 16'd 7832;
    assign memory[3739] = 16'd 7854;
    assign memory[3740] = 16'd 7875;
    assign memory[3741] = 16'd 7897;
    assign memory[3742] = 16'd 7918;
    assign memory[3743] = 16'd 7940;
    assign memory[3744] = 16'd 7961;
    assign memory[3745] = 16'd 7983;
    assign memory[3746] = 16'd 8005;
    assign memory[3747] = 16'd 8026;
    assign memory[3748] = 16'd 8048;
    assign memory[3749] = 16'd 8069;
    assign memory[3750] = 16'd 8091;
    assign memory[3751] = 16'd 8113;
    assign memory[3752] = 16'd 8135;
    assign memory[3753] = 16'd 8156;
    assign memory[3754] = 16'd 8178;
    assign memory[3755] = 16'd 8200;
    assign memory[3756] = 16'd 8222;
    assign memory[3757] = 16'd 8243;
    assign memory[3758] = 16'd 8265;
    assign memory[3759] = 16'd 8287;
    assign memory[3760] = 16'd 8309;
    assign memory[3761] = 16'd 8331;
    assign memory[3762] = 16'd 8353;
    assign memory[3763] = 16'd 8375;
    assign memory[3764] = 16'd 8396;
    assign memory[3765] = 16'd 8418;
    assign memory[3766] = 16'd 8440;
    assign memory[3767] = 16'd 8462;
    assign memory[3768] = 16'd 8484;
    assign memory[3769] = 16'd 8506;
    assign memory[3770] = 16'd 8528;
    assign memory[3771] = 16'd 8551;
    assign memory[3772] = 16'd 8573;
    assign memory[3773] = 16'd 8595;
    assign memory[3774] = 16'd 8617;
    assign memory[3775] = 16'd 8639;
    assign memory[3776] = 16'd 8661;
    assign memory[3777] = 16'd 8683;
    assign memory[3778] = 16'd 8706;
    assign memory[3779] = 16'd 8728;
    assign memory[3780] = 16'd 8750;
    assign memory[3781] = 16'd 8772;
    assign memory[3782] = 16'd 8794;
    assign memory[3783] = 16'd 8817;
    assign memory[3784] = 16'd 8839;
    assign memory[3785] = 16'd 8861;
    assign memory[3786] = 16'd 8884;
    assign memory[3787] = 16'd 8906;
    assign memory[3788] = 16'd 8928;
    assign memory[3789] = 16'd 8951;
    assign memory[3790] = 16'd 8973;
    assign memory[3791] = 16'd 8996;
    assign memory[3792] = 16'd 9018;
    assign memory[3793] = 16'd 9041;
    assign memory[3794] = 16'd 9063;
    assign memory[3795] = 16'd 9085;
    assign memory[3796] = 16'd 9108;
    assign memory[3797] = 16'd 9131;
    assign memory[3798] = 16'd 9153;
    assign memory[3799] = 16'd 9176;
    assign memory[3800] = 16'd 9198;
    assign memory[3801] = 16'd 9221;
    assign memory[3802] = 16'd 9243;
    assign memory[3803] = 16'd 9266;
    assign memory[3804] = 16'd 9289;
    assign memory[3805] = 16'd 9311;
    assign memory[3806] = 16'd 9334;
    assign memory[3807] = 16'd 9357;
    assign memory[3808] = 16'd 9379;
    assign memory[3809] = 16'd 9402;
    assign memory[3810] = 16'd 9425;
    assign memory[3811] = 16'd 9448;
    assign memory[3812] = 16'd 9470;
    assign memory[3813] = 16'd 9493;
    assign memory[3814] = 16'd 9516;
    assign memory[3815] = 16'd 9539;
    assign memory[3816] = 16'd 9562;
    assign memory[3817] = 16'd 9585;
    assign memory[3818] = 16'd 9607;
    assign memory[3819] = 16'd 9630;
    assign memory[3820] = 16'd 9653;
    assign memory[3821] = 16'd 9676;
    assign memory[3822] = 16'd 9699;
    assign memory[3823] = 16'd 9722;
    assign memory[3824] = 16'd 9745;
    assign memory[3825] = 16'd 9768;
    assign memory[3826] = 16'd 9791;
    assign memory[3827] = 16'd 9814;
    assign memory[3828] = 16'd 9837;
    assign memory[3829] = 16'd 9860;
    assign memory[3830] = 16'd 9883;
    assign memory[3831] = 16'd 9906;
    assign memory[3832] = 16'd 9929;
    assign memory[3833] = 16'd 9952;
    assign memory[3834] = 16'd 9976;
    assign memory[3835] = 16'd 9999;
    assign memory[3836] = 16'd10022;
    assign memory[3837] = 16'd10045;
    assign memory[3838] = 16'd10068;
    assign memory[3839] = 16'd10091;
    assign memory[3840] = 16'd10115;
    assign memory[3841] = 16'd10138;
    assign memory[3842] = 16'd10161;
    assign memory[3843] = 16'd10184;
    assign memory[3844] = 16'd10208;
    assign memory[3845] = 16'd10231;
    assign memory[3846] = 16'd10254;
    assign memory[3847] = 16'd10278;
    assign memory[3848] = 16'd10301;
    assign memory[3849] = 16'd10324;
    assign memory[3850] = 16'd10348;
    assign memory[3851] = 16'd10371;
    assign memory[3852] = 16'd10394;
    assign memory[3853] = 16'd10418;
    assign memory[3854] = 16'd10441;
    assign memory[3855] = 16'd10465;
    assign memory[3856] = 16'd10488;
    assign memory[3857] = 16'd10511;
    assign memory[3858] = 16'd10535;
    assign memory[3859] = 16'd10558;
    assign memory[3860] = 16'd10582;
    assign memory[3861] = 16'd10605;
    assign memory[3862] = 16'd10629;
    assign memory[3863] = 16'd10652;
    assign memory[3864] = 16'd10676;
    assign memory[3865] = 16'd10700;
    assign memory[3866] = 16'd10723;
    assign memory[3867] = 16'd10747;
    assign memory[3868] = 16'd10770;
    assign memory[3869] = 16'd10794;
    assign memory[3870] = 16'd10818;
    assign memory[3871] = 16'd10841;
    assign memory[3872] = 16'd10865;
    assign memory[3873] = 16'd10889;
    assign memory[3874] = 16'd10912;
    assign memory[3875] = 16'd10936;
    assign memory[3876] = 16'd10960;
    assign memory[3877] = 16'd10983;
    assign memory[3878] = 16'd11007;
    assign memory[3879] = 16'd11031;
    assign memory[3880] = 16'd11055;
    assign memory[3881] = 16'd11078;
    assign memory[3882] = 16'd11102;
    assign memory[3883] = 16'd11126;
    assign memory[3884] = 16'd11150;
    assign memory[3885] = 16'd11174;
    assign memory[3886] = 16'd11197;
    assign memory[3887] = 16'd11221;
    assign memory[3888] = 16'd11245;
    assign memory[3889] = 16'd11269;
    assign memory[3890] = 16'd11293;
    assign memory[3891] = 16'd11317;
    assign memory[3892] = 16'd11341;
    assign memory[3893] = 16'd11365;
    assign memory[3894] = 16'd11389;
    assign memory[3895] = 16'd11412;
    assign memory[3896] = 16'd11436;
    assign memory[3897] = 16'd11460;
    assign memory[3898] = 16'd11484;
    assign memory[3899] = 16'd11508;
    assign memory[3900] = 16'd11532;
    assign memory[3901] = 16'd11556;
    assign memory[3902] = 16'd11580;
    assign memory[3903] = 16'd11604;
    assign memory[3904] = 16'd11628;
    assign memory[3905] = 16'd11653;
    assign memory[3906] = 16'd11677;
    assign memory[3907] = 16'd11701;
    assign memory[3908] = 16'd11725;
    assign memory[3909] = 16'd11749;
    assign memory[3910] = 16'd11773;
    assign memory[3911] = 16'd11797;
    assign memory[3912] = 16'd11821;
    assign memory[3913] = 16'd11845;
    assign memory[3914] = 16'd11870;
    assign memory[3915] = 16'd11894;
    assign memory[3916] = 16'd11918;
    assign memory[3917] = 16'd11942;
    assign memory[3918] = 16'd11966;
    assign memory[3919] = 16'd11990;
    assign memory[3920] = 16'd12015;
    assign memory[3921] = 16'd12039;
    assign memory[3922] = 16'd12063;
    assign memory[3923] = 16'd12087;
    assign memory[3924] = 16'd12112;
    assign memory[3925] = 16'd12136;
    assign memory[3926] = 16'd12160;
    assign memory[3927] = 16'd12184;
    assign memory[3928] = 16'd12209;
    assign memory[3929] = 16'd12233;
    assign memory[3930] = 16'd12257;
    assign memory[3931] = 16'd12282;
    assign memory[3932] = 16'd12306;
    assign memory[3933] = 16'd12330;
    assign memory[3934] = 16'd12355;
    assign memory[3935] = 16'd12379;
    assign memory[3936] = 16'd12404;
    assign memory[3937] = 16'd12428;
    assign memory[3938] = 16'd12452;
    assign memory[3939] = 16'd12477;
    assign memory[3940] = 16'd12501;
    assign memory[3941] = 16'd12526;
    assign memory[3942] = 16'd12550;
    assign memory[3943] = 16'd12574;
    assign memory[3944] = 16'd12599;
    assign memory[3945] = 16'd12623;
    assign memory[3946] = 16'd12648;
    assign memory[3947] = 16'd12672;
    assign memory[3948] = 16'd12697;
    assign memory[3949] = 16'd12721;
    assign memory[3950] = 16'd12746;
    assign memory[3951] = 16'd12770;
    assign memory[3952] = 16'd12795;
    assign memory[3953] = 16'd12819;
    assign memory[3954] = 16'd12844;
    assign memory[3955] = 16'd12868;
    assign memory[3956] = 16'd12893;
    assign memory[3957] = 16'd12917;
    assign memory[3958] = 16'd12942;
    assign memory[3959] = 16'd12967;
    assign memory[3960] = 16'd12991;
    assign memory[3961] = 16'd13016;
    assign memory[3962] = 16'd13040;
    assign memory[3963] = 16'd13065;
    assign memory[3964] = 16'd13090;
    assign memory[3965] = 16'd13114;
    assign memory[3966] = 16'd13139;
    assign memory[3967] = 16'd13163;
    assign memory[3968] = 16'd13188;
    assign memory[3969] = 16'd13213;
    assign memory[3970] = 16'd13237;
    assign memory[3971] = 16'd13262;
    assign memory[3972] = 16'd13287;
    assign memory[3973] = 16'd13311;
    assign memory[3974] = 16'd13336;
    assign memory[3975] = 16'd13361;
    assign memory[3976] = 16'd13386;
    assign memory[3977] = 16'd13410;
    assign memory[3978] = 16'd13435;
    assign memory[3979] = 16'd13460;
    assign memory[3980] = 16'd13484;
    assign memory[3981] = 16'd13509;
    assign memory[3982] = 16'd13534;
    assign memory[3983] = 16'd13559;
    assign memory[3984] = 16'd13583;
    assign memory[3985] = 16'd13608;
    assign memory[3986] = 16'd13633;
    assign memory[3987] = 16'd13658;
    assign memory[3988] = 16'd13683;
    assign memory[3989] = 16'd13707;
    assign memory[3990] = 16'd13732;
    assign memory[3991] = 16'd13757;
    assign memory[3992] = 16'd13782;
    assign memory[3993] = 16'd13807;
    assign memory[3994] = 16'd13831;
    assign memory[3995] = 16'd13856;
    assign memory[3996] = 16'd13881;
    assign memory[3997] = 16'd13906;
    assign memory[3998] = 16'd13931;
    assign memory[3999] = 16'd13956;
    assign memory[4000] = 16'd13980;
    assign memory[4001] = 16'd14005;
    assign memory[4002] = 16'd14030;
    assign memory[4003] = 16'd14055;
    assign memory[4004] = 16'd14080;
    assign memory[4005] = 16'd14105;
    assign memory[4006] = 16'd14130;
    assign memory[4007] = 16'd14155;
    assign memory[4008] = 16'd14180;
    assign memory[4009] = 16'd14204;
    assign memory[4010] = 16'd14229;
    assign memory[4011] = 16'd14254;
    assign memory[4012] = 16'd14279;
    assign memory[4013] = 16'd14304;
    assign memory[4014] = 16'd14329;
    assign memory[4015] = 16'd14354;
    assign memory[4016] = 16'd14379;
    assign memory[4017] = 16'd14404;
    assign memory[4018] = 16'd14429;
    assign memory[4019] = 16'd14454;
    assign memory[4020] = 16'd14479;
    assign memory[4021] = 16'd14504;
    assign memory[4022] = 16'd14529;
    assign memory[4023] = 16'd14554;
    assign memory[4024] = 16'd14579;
    assign memory[4025] = 16'd14604;
    assign memory[4026] = 16'd14629;
    assign memory[4027] = 16'd14654;
    assign memory[4028] = 16'd14679;
    assign memory[4029] = 16'd14704;
    assign memory[4030] = 16'd14729;
    assign memory[4031] = 16'd14754;
    assign memory[4032] = 16'd14779;
    assign memory[4033] = 16'd14804;
    assign memory[4034] = 16'd14829;
    assign memory[4035] = 16'd14854;
    assign memory[4036] = 16'd14879;
    assign memory[4037] = 16'd14904;
    assign memory[4038] = 16'd14929;
    assign memory[4039] = 16'd14954;
    assign memory[4040] = 16'd14979;
    assign memory[4041] = 16'd15004;
    assign memory[4042] = 16'd15029;
    assign memory[4043] = 16'd15054;
    assign memory[4044] = 16'd15079;
    assign memory[4045] = 16'd15104;
    assign memory[4046] = 16'd15129;
    assign memory[4047] = 16'd15154;
    assign memory[4048] = 16'd15179;
    assign memory[4049] = 16'd15204;
    assign memory[4050] = 16'd15229;
    assign memory[4051] = 16'd15254;
    assign memory[4052] = 16'd15279;
    assign memory[4053] = 16'd15305;
    assign memory[4054] = 16'd15330;
    assign memory[4055] = 16'd15355;
    assign memory[4056] = 16'd15380;
    assign memory[4057] = 16'd15405;
    assign memory[4058] = 16'd15430;
    assign memory[4059] = 16'd15455;
    assign memory[4060] = 16'd15480;
    assign memory[4061] = 16'd15505;
    assign memory[4062] = 16'd15530;
    assign memory[4063] = 16'd15555;
    assign memory[4064] = 16'd15581;
    assign memory[4065] = 16'd15606;
    assign memory[4066] = 16'd15631;
    assign memory[4067] = 16'd15656;
    assign memory[4068] = 16'd15681;
    assign memory[4069] = 16'd15706;
    assign memory[4070] = 16'd15731;
    assign memory[4071] = 16'd15756;
    assign memory[4072] = 16'd15781;
    assign memory[4073] = 16'd15807;
    assign memory[4074] = 16'd15832;
    assign memory[4075] = 16'd15857;
    assign memory[4076] = 16'd15882;
    assign memory[4077] = 16'd15907;
    assign memory[4078] = 16'd15932;
    assign memory[4079] = 16'd15957;
    assign memory[4080] = 16'd15982;
    assign memory[4081] = 16'd16008;
    assign memory[4082] = 16'd16033;
    assign memory[4083] = 16'd16058;
    assign memory[4084] = 16'd16083;
    assign memory[4085] = 16'd16108;
    assign memory[4086] = 16'd16133;
    assign memory[4087] = 16'd16158;
    assign memory[4088] = 16'd16183;
    assign memory[4089] = 16'd16209;
    assign memory[4090] = 16'd16234;
    assign memory[4091] = 16'd16259;
    assign memory[4092] = 16'd16284;
    assign memory[4093] = 16'd16309;
    assign memory[4094] = 16'd16334;
    assign memory[4095] = 16'd16359;

endmodule
