module lead_rom (
    input clk,
	output reg [15:0] dout,
	input [11:0] addr
    );
	
	wire [15:0] memory [543:0];

	always @(posedge clk) begin
        if (addr < 12'd544) begin
            dout = memory[addr];
        end else if (addr < 12'd3584) begin
            dout = 16'd32767;
        end else begin
            dout = 16'd0;
        end
    end
    
    assign memory[0   ] = 16'd0    ;
    assign memory[1   ] = 16'd543  ;
    assign memory[2   ] = 16'd1078 ;
    assign memory[3   ] = 16'd1605 ;
    assign memory[4   ] = 16'd2123 ;
    assign memory[5   ] = 16'd2634 ;
    assign memory[6   ] = 16'd3136 ;
    assign memory[7   ] = 16'd3631 ;
    assign memory[8   ] = 16'd4118 ;
    assign memory[9   ] = 16'd4598 ;
    assign memory[10  ] = 16'd5070 ;
    assign memory[11  ] = 16'd5534 ;
    assign memory[12  ] = 16'd5991 ;
    assign memory[13  ] = 16'd6441 ;
    assign memory[14  ] = 16'd6884 ;
    assign memory[15  ] = 16'd7320 ;
    assign memory[16  ] = 16'd7748 ;
    assign memory[17  ] = 16'd8170 ;
    assign memory[18  ] = 16'd8585 ;
    assign memory[19  ] = 16'd8994 ;
    assign memory[20  ] = 16'd9395 ;
    assign memory[21  ] = 16'd9791 ;
    assign memory[22  ] = 16'd10179;
    assign memory[23  ] = 16'd10562;
    assign memory[24  ] = 16'd10938;
    assign memory[25  ] = 16'd11308;
    assign memory[26  ] = 16'd11672;
    assign memory[27  ] = 16'd12030;
    assign memory[28  ] = 16'd12382;
    assign memory[29  ] = 16'd12729;
    assign memory[30  ] = 16'd13069;
    assign memory[31  ] = 16'd13404;
    assign memory[32  ] = 16'd13733;
    assign memory[33  ] = 16'd14057;
    assign memory[34  ] = 16'd14375;
    assign memory[35  ] = 16'd14688;
    assign memory[36  ] = 16'd14996;
    assign memory[37  ] = 16'd15298;
    assign memory[38  ] = 16'd15595;
    assign memory[39  ] = 16'd15887;
    assign memory[40  ] = 16'd16175;
    assign memory[41  ] = 16'd16457;
    assign memory[42  ] = 16'd16734;
    assign memory[43  ] = 16'd17007;
    assign memory[44  ] = 16'd17275;
    assign memory[45  ] = 16'd17538;
    assign memory[46  ] = 16'd17797;
    assign memory[47  ] = 16'd18051;
    assign memory[48  ] = 16'd18301;
    assign memory[49  ] = 16'd18546;
    assign memory[50  ] = 16'd18788;
    assign memory[51  ] = 16'd19024;
    assign memory[52  ] = 16'd19257;
    assign memory[53  ] = 16'd19486;
    assign memory[54  ] = 16'd19710;
    assign memory[55  ] = 16'd19931;
    assign memory[56  ] = 16'd20147;
    assign memory[57  ] = 16'd20360;
    assign memory[58  ] = 16'd20569;
    assign memory[59  ] = 16'd20774;
    assign memory[60  ] = 16'd20975;
    assign memory[61  ] = 16'd21173;
    assign memory[62  ] = 16'd21367;
    assign memory[63  ] = 16'd21558;
    assign memory[64  ] = 16'd21745;
    assign memory[65  ] = 16'd21929;
    assign memory[66  ] = 16'd22109;
    assign memory[67  ] = 16'd22286;
    assign memory[68  ] = 16'd22460;
    assign memory[69  ] = 16'd22631;
    assign memory[70  ] = 16'd22798;
    assign memory[71  ] = 16'd22963;
    assign memory[72  ] = 16'd23124;
    assign memory[73  ] = 16'd23283;
    assign memory[74  ] = 16'd23438;
    assign memory[75  ] = 16'd23590;
    assign memory[76  ] = 16'd23740;
    assign memory[77  ] = 16'd23887;
    assign memory[78  ] = 16'd24031;
    assign memory[79  ] = 16'd24172;
    assign memory[80  ] = 16'd24311;
    assign memory[81  ] = 16'd24447;
    assign memory[82  ] = 16'd24580;
    assign memory[83  ] = 16'd24711;
    assign memory[84  ] = 16'd24840;
    assign memory[85  ] = 16'd24965;
    assign memory[86  ] = 16'd25089;
    assign memory[87  ] = 16'd25210;
    assign memory[88  ] = 16'd25329;
    assign memory[89  ] = 16'd25445;
    assign memory[90  ] = 16'd25560;
    assign memory[91  ] = 16'd25672;
    assign memory[92  ] = 16'd25782;
    assign memory[93  ] = 16'd25890;
    assign memory[94  ] = 16'd25995;
    assign memory[95  ] = 16'd26099;
    assign memory[96  ] = 16'd26200;
    assign memory[97  ] = 16'd26300;
    assign memory[98  ] = 16'd26398;
    assign memory[99  ] = 16'd26493;
    assign memory[100 ] = 16'd26587;
    assign memory[101 ] = 16'd26679;
    assign memory[102 ] = 16'd26770;
    assign memory[103 ] = 16'd26858;
    assign memory[104 ] = 16'd26945;
    assign memory[105 ] = 16'd27030;
    assign memory[106 ] = 16'd27113;
    assign memory[107 ] = 16'd27195;
    assign memory[108 ] = 16'd27275;
    assign memory[109 ] = 16'd27353;
    assign memory[110 ] = 16'd27430;
    assign memory[111 ] = 16'd27505;
    assign memory[112 ] = 16'd27579;
    assign memory[113 ] = 16'd27651;
    assign memory[114 ] = 16'd27722;
    assign memory[115 ] = 16'd27792;
    assign memory[116 ] = 16'd27860;
    assign memory[117 ] = 16'd27927;
    assign memory[118 ] = 16'd27992;
    assign memory[119 ] = 16'd28056;
    assign memory[120 ] = 16'd28119;
    assign memory[121 ] = 16'd28181;
    assign memory[122 ] = 16'd28241;
    assign memory[123 ] = 16'd28300;
    assign memory[124 ] = 16'd28358;
    assign memory[125 ] = 16'd28415;
    assign memory[126 ] = 16'd28471;
    assign memory[127 ] = 16'd28526;
    assign memory[128 ] = 16'd28579;
    assign memory[129 ] = 16'd28631;
    assign memory[130 ] = 16'd28683;
    assign memory[131 ] = 16'd28733;
    assign memory[132 ] = 16'd28783;
    assign memory[133 ] = 16'd28831;
    assign memory[134 ] = 16'd28878;
    assign memory[135 ] = 16'd28925;
    assign memory[136 ] = 16'd28970;
    assign memory[137 ] = 16'd29015;
    assign memory[138 ] = 16'd29059;
    assign memory[139 ] = 16'd29102;
    assign memory[140 ] = 16'd29144;
    assign memory[141 ] = 16'd29185;
    assign memory[142 ] = 16'd29226;
    assign memory[143 ] = 16'd29265;
    assign memory[144 ] = 16'd29304;
    assign memory[145 ] = 16'd29342;
    assign memory[146 ] = 16'd29380;
    assign memory[147 ] = 16'd29417;
    assign memory[148 ] = 16'd29453;
    assign memory[149 ] = 16'd29488;
    assign memory[150 ] = 16'd29522;
    assign memory[151 ] = 16'd29556;
    assign memory[152 ] = 16'd29590;
    assign memory[153 ] = 16'd29622;
    assign memory[154 ] = 16'd29655;
    assign memory[155 ] = 16'd29686;
    assign memory[156 ] = 16'd29717;
    assign memory[157 ] = 16'd29747;
    assign memory[158 ] = 16'd29777;
    assign memory[159 ] = 16'd29806;
    assign memory[160 ] = 16'd29835;
    assign memory[161 ] = 16'd29863;
    assign memory[162 ] = 16'd29891;
    assign memory[163 ] = 16'd29918;
    assign memory[164 ] = 16'd29944;
    assign memory[165 ] = 16'd29971;
    assign memory[166 ] = 16'd29996;
    assign memory[167 ] = 16'd30022;
    assign memory[168 ] = 16'd30046;
    assign memory[169 ] = 16'd30071;
    assign memory[170 ] = 16'd30095;
    assign memory[171 ] = 16'd30118;
    assign memory[172 ] = 16'd30142;
    assign memory[173 ] = 16'd30164;
    assign memory[174 ] = 16'd30187;
    assign memory[175 ] = 16'd30209;
    assign memory[176 ] = 16'd30231;
    assign memory[177 ] = 16'd30252;
    assign memory[178 ] = 16'd30273;
    assign memory[179 ] = 16'd30293;
    assign memory[180 ] = 16'd30314;
    assign memory[181 ] = 16'd30334;
    assign memory[182 ] = 16'd30353;
    assign memory[183 ] = 16'd30373;
    assign memory[184 ] = 16'd30392;
    assign memory[185 ] = 16'd30411;
    assign memory[186 ] = 16'd30429;
    assign memory[187 ] = 16'd30447;
    assign memory[188 ] = 16'd30465;
    assign memory[189 ] = 16'd30483;
    assign memory[190 ] = 16'd30500;
    assign memory[191 ] = 16'd30517;
    assign memory[192 ] = 16'd30534;
    assign memory[193 ] = 16'd30551;
    assign memory[194 ] = 16'd30568;
    assign memory[195 ] = 16'd30584;
    assign memory[196 ] = 16'd30600;
    assign memory[197 ] = 16'd30616;
    assign memory[198 ] = 16'd30631;
    assign memory[199 ] = 16'd30646;
    assign memory[200 ] = 16'd30662;
    assign memory[201 ] = 16'd30677;
    assign memory[202 ] = 16'd30691;
    assign memory[203 ] = 16'd30706;
    assign memory[204 ] = 16'd30720;
    assign memory[205 ] = 16'd30735;
    assign memory[206 ] = 16'd30749;
    assign memory[207 ] = 16'd30763;
    assign memory[208 ] = 16'd30776;
    assign memory[209 ] = 16'd30790;
    assign memory[210 ] = 16'd30803;
    assign memory[211 ] = 16'd30816;
    assign memory[212 ] = 16'd30829;
    assign memory[213 ] = 16'd30842;
    assign memory[214 ] = 16'd30855;
    assign memory[215 ] = 16'd30868;
    assign memory[216 ] = 16'd30880;
    assign memory[217 ] = 16'd30893;
    assign memory[218 ] = 16'd30905;
    assign memory[219 ] = 16'd30917;
    assign memory[220 ] = 16'd30929;
    assign memory[221 ] = 16'd30941;
    assign memory[222 ] = 16'd30952;
    assign memory[223 ] = 16'd30964;
    assign memory[224 ] = 16'd30975;
    assign memory[225 ] = 16'd30987;
    assign memory[226 ] = 16'd30998;
    assign memory[227 ] = 16'd31009;
    assign memory[228 ] = 16'd31020;
    assign memory[229 ] = 16'd31031;
    assign memory[230 ] = 16'd31042;
    assign memory[231 ] = 16'd31052;
    assign memory[232 ] = 16'd31063;
    assign memory[233 ] = 16'd31073;
    assign memory[234 ] = 16'd31084;
    assign memory[235 ] = 16'd31094;
    assign memory[236 ] = 16'd31104;
    assign memory[237 ] = 16'd31114;
    assign memory[238 ] = 16'd31124;
    assign memory[239 ] = 16'd31134;
    assign memory[240 ] = 16'd31143;
    assign memory[241 ] = 16'd31153;
    assign memory[242 ] = 16'd31163;
    assign memory[243 ] = 16'd31172;
    assign memory[244 ] = 16'd31181;
    assign memory[245 ] = 16'd31191;
    assign memory[246 ] = 16'd31200;
    assign memory[247 ] = 16'd31209;
    assign memory[248 ] = 16'd31218;
    assign memory[249 ] = 16'd31227;
    assign memory[250 ] = 16'd31235;
    assign memory[251 ] = 16'd31244;
    assign memory[252 ] = 16'd31253;
    assign memory[253 ] = 16'd31261;
    assign memory[254 ] = 16'd31269;
    assign memory[255 ] = 16'd31278;
    assign memory[256 ] = 16'd31286;
    assign memory[257 ] = 16'd31294;
    assign memory[258 ] = 16'd31302;
    assign memory[259 ] = 16'd31310;
    assign memory[260 ] = 16'd31318;
    assign memory[261 ] = 16'd31326;
    assign memory[262 ] = 16'd31334;
    assign memory[263 ] = 16'd31341;
    assign memory[264 ] = 16'd31349;
    assign memory[265 ] = 16'd31356;
    assign memory[266 ] = 16'd31364;
    assign memory[267 ] = 16'd31371;
    assign memory[268 ] = 16'd31378;
    assign memory[269 ] = 16'd31385;
    assign memory[270 ] = 16'd31392;
    assign memory[271 ] = 16'd31399;
    assign memory[272 ] = 16'd31406;
    assign memory[273 ] = 16'd31413;
    assign memory[274 ] = 16'd31419;
    assign memory[275 ] = 16'd31426;
    assign memory[276 ] = 16'd31432;
    assign memory[277 ] = 16'd31439;
    assign memory[278 ] = 16'd31445;
    assign memory[279 ] = 16'd31451;
    assign memory[280 ] = 16'd31458;
    assign memory[281 ] = 16'd31464;
    assign memory[282 ] = 16'd31470;
    assign memory[283 ] = 16'd31475;
    assign memory[284 ] = 16'd31481;
    assign memory[285 ] = 16'd31487;
    assign memory[286 ] = 16'd31493;
    assign memory[287 ] = 16'd31498;
    assign memory[288 ] = 16'd31504;
    assign memory[289 ] = 16'd31509;
    assign memory[290 ] = 16'd31514;
    assign memory[291 ] = 16'd31519;
    assign memory[292 ] = 16'd31525;
    assign memory[293 ] = 16'd31530;
    assign memory[294 ] = 16'd31534;
    assign memory[295 ] = 16'd31539;
    assign memory[296 ] = 16'd31544;
    assign memory[297 ] = 16'd31549;
    assign memory[298 ] = 16'd31553;
    assign memory[299 ] = 16'd31558;
    assign memory[300 ] = 16'd31562;
    assign memory[301 ] = 16'd31567;
    assign memory[302 ] = 16'd31571;
    assign memory[303 ] = 16'd31575;
    assign memory[304 ] = 16'd31579;
    assign memory[305 ] = 16'd31583;
    assign memory[306 ] = 16'd31587;
    assign memory[307 ] = 16'd31591;
    assign memory[308 ] = 16'd31595;
    assign memory[309 ] = 16'd31598;
    assign memory[310 ] = 16'd31602;
    assign memory[311 ] = 16'd31605;
    assign memory[312 ] = 16'd31609;
    assign memory[313 ] = 16'd31612;
    assign memory[314 ] = 16'd31616;
    assign memory[315 ] = 16'd31619;
    assign memory[316 ] = 16'd31622;
    assign memory[317 ] = 16'd31625;
    assign memory[318 ] = 16'd31628;
    assign memory[319 ] = 16'd31631;
    assign memory[320 ] = 16'd31634;
    assign memory[321 ] = 16'd31636;
    assign memory[322 ] = 16'd31639;
    assign memory[323 ] = 16'd31642;
    assign memory[324 ] = 16'd31644;
    assign memory[325 ] = 16'd31646;
    assign memory[326 ] = 16'd31649;
    assign memory[327 ] = 16'd31651;
    assign memory[328 ] = 16'd31653;
    assign memory[329 ] = 16'd31656;
    assign memory[330 ] = 16'd31658;
    assign memory[331 ] = 16'd31660;
    assign memory[332 ] = 16'd31662;
    assign memory[333 ] = 16'd31664;
    assign memory[334 ] = 16'd31665;
    assign memory[335 ] = 16'd31667;
    assign memory[336 ] = 16'd31669;
    assign memory[337 ] = 16'd31670;
    assign memory[338 ] = 16'd31672;
    assign memory[339 ] = 16'd31674;
    assign memory[340 ] = 16'd31675;
    assign memory[341 ] = 16'd31676;
    assign memory[342 ] = 16'd31678;
    assign memory[343 ] = 16'd31679;
    assign memory[344 ] = 16'd31680;
    assign memory[345 ] = 16'd31682;
    assign memory[346 ] = 16'd31683;
    assign memory[347 ] = 16'd31684;
    assign memory[348 ] = 16'd31685;
    assign memory[349 ] = 16'd31686;
    assign memory[350 ] = 16'd31687;
    assign memory[351 ] = 16'd31688;
    assign memory[352 ] = 16'd31689;
    assign memory[353 ] = 16'd31690;
    assign memory[354 ] = 16'd31691;
    assign memory[355 ] = 16'd31692;
    assign memory[356 ] = 16'd31692;
    assign memory[357 ] = 16'd31693;
    assign memory[358 ] = 16'd31694;
    assign memory[359 ] = 16'd31694;
    assign memory[360 ] = 16'd31695;
    assign memory[361 ] = 16'd31696;
    assign memory[362 ] = 16'd31696;
    assign memory[363 ] = 16'd31697;
    assign memory[364 ] = 16'd31698;
    assign memory[365 ] = 16'd31698;
    assign memory[366 ] = 16'd31699;
    assign memory[367 ] = 16'd31699;
    assign memory[368 ] = 16'd31700;
    assign memory[369 ] = 16'd31700;
    assign memory[370 ] = 16'd31701;
    assign memory[371 ] = 16'd31702;
    assign memory[372 ] = 16'd31702;
    assign memory[373 ] = 16'd31703;
    assign memory[374 ] = 16'd31703;
    assign memory[375 ] = 16'd31704;
    assign memory[376 ] = 16'd31704;
    assign memory[377 ] = 16'd31705;
    assign memory[378 ] = 16'd31705;
    assign memory[379 ] = 16'd31706;
    assign memory[380 ] = 16'd31707;
    assign memory[381 ] = 16'd31707;
    assign memory[382 ] = 16'd31708;
    assign memory[383 ] = 16'd31709;
    assign memory[384 ] = 16'd31709;
    assign memory[385 ] = 16'd31710;
    assign memory[386 ] = 16'd31711;
    assign memory[387 ] = 16'd31712;
    assign memory[388 ] = 16'd31713;
    assign memory[389 ] = 16'd31713;
    assign memory[390 ] = 16'd31714;
    assign memory[391 ] = 16'd31715;
    assign memory[392 ] = 16'd31716;
    assign memory[393 ] = 16'd31717;
    assign memory[394 ] = 16'd31718;
    assign memory[395 ] = 16'd31720;
    assign memory[396 ] = 16'd31721;
    assign memory[397 ] = 16'd31722;
    assign memory[398 ] = 16'd31723;
    assign memory[399 ] = 16'd31725;
    assign memory[400 ] = 16'd31726;
    assign memory[401 ] = 16'd31728;
    assign memory[402 ] = 16'd31729;
    assign memory[403 ] = 16'd31731;
    assign memory[404 ] = 16'd31733;
    assign memory[405 ] = 16'd31735;
    assign memory[406 ] = 16'd31736;
    assign memory[407 ] = 16'd31738;
    assign memory[408 ] = 16'd31741;
    assign memory[409 ] = 16'd31743;
    assign memory[410 ] = 16'd31745;
    assign memory[411 ] = 16'd31747;
    assign memory[412 ] = 16'd31750;
    assign memory[413 ] = 16'd31752;
    assign memory[414 ] = 16'd31755;
    assign memory[415 ] = 16'd31757;
    assign memory[416 ] = 16'd31760;
    assign memory[417 ] = 16'd31763;
    assign memory[418 ] = 16'd31766;
    assign memory[419 ] = 16'd31769;
    assign memory[420 ] = 16'd31772;
    assign memory[421 ] = 16'd31776;
    assign memory[422 ] = 16'd31779;
    assign memory[423 ] = 16'd31783;
    assign memory[424 ] = 16'd31786;
    assign memory[425 ] = 16'd31790;
    assign memory[426 ] = 16'd31794;
    assign memory[427 ] = 16'd31798;
    assign memory[428 ] = 16'd31802;
    assign memory[429 ] = 16'd31806;
    assign memory[430 ] = 16'd31811;
    assign memory[431 ] = 16'd31815;
    assign memory[432 ] = 16'd31820;
    assign memory[433 ] = 16'd31825;
    assign memory[434 ] = 16'd31829;
    assign memory[435 ] = 16'd31834;
    assign memory[436 ] = 16'd31840;
    assign memory[437 ] = 16'd31845;
    assign memory[438 ] = 16'd31850;
    assign memory[439 ] = 16'd31856;
    assign memory[440 ] = 16'd31862;
    assign memory[441 ] = 16'd31867;
    assign memory[442 ] = 16'd31873;
    assign memory[443 ] = 16'd31879;
    assign memory[444 ] = 16'd31886;
    assign memory[445 ] = 16'd31892;
    assign memory[446 ] = 16'd31899;
    assign memory[447 ] = 16'd31905;
    assign memory[448 ] = 16'd31912;
    assign memory[449 ] = 16'd31919;
    assign memory[450 ] = 16'd31926;
    assign memory[451 ] = 16'd31933;
    assign memory[452 ] = 16'd31941;
    assign memory[453 ] = 16'd31948;
    assign memory[454 ] = 16'd31956;
    assign memory[455 ] = 16'd31963;
    assign memory[456 ] = 16'd31971;
    assign memory[457 ] = 16'd31979;
    assign memory[458 ] = 16'd31988;
    assign memory[459 ] = 16'd31996;
    assign memory[460 ] = 16'd32004;
    assign memory[461 ] = 16'd32013;
    assign memory[462 ] = 16'd32022;
    assign memory[463 ] = 16'd32031;
    assign memory[464 ] = 16'd32040;
    assign memory[465 ] = 16'd32049;
    assign memory[466 ] = 16'd32058;
    assign memory[467 ] = 16'd32067;
    assign memory[468 ] = 16'd32077;
    assign memory[469 ] = 16'd32087;
    assign memory[470 ] = 16'd32096;
    assign memory[471 ] = 16'd32106;
    assign memory[472 ] = 16'd32116;
    assign memory[473 ] = 16'd32126;
    assign memory[474 ] = 16'd32137;
    assign memory[475 ] = 16'd32147;
    assign memory[476 ] = 16'd32157;
    assign memory[477 ] = 16'd32168;
    assign memory[478 ] = 16'd32178;
    assign memory[479 ] = 16'd32189;
    assign memory[480 ] = 16'd32200;
    assign memory[481 ] = 16'd32211;
    assign memory[482 ] = 16'd32222;
    assign memory[483 ] = 16'd32233;
    assign memory[484 ] = 16'd32244;
    assign memory[485 ] = 16'd32255;
    assign memory[486 ] = 16'd32267;
    assign memory[487 ] = 16'd32278;
    assign memory[488 ] = 16'd32289;
    assign memory[489 ] = 16'd32301;
    assign memory[490 ] = 16'd32312;
    assign memory[491 ] = 16'd32324;
    assign memory[492 ] = 16'd32335;
    assign memory[493 ] = 16'd32347;
    assign memory[494 ] = 16'd32359;
    assign memory[495 ] = 16'd32370;
    assign memory[496 ] = 16'd32382;
    assign memory[497 ] = 16'd32394;
    assign memory[498 ] = 16'd32405;
    assign memory[499 ] = 16'd32417;
    assign memory[500 ] = 16'd32429;
    assign memory[501 ] = 16'd32440;
    assign memory[502 ] = 16'd32452;
    assign memory[503 ] = 16'd32463;
    assign memory[504 ] = 16'd32475;
    assign memory[505 ] = 16'd32486;
    assign memory[506 ] = 16'd32498;
    assign memory[507 ] = 16'd32509;
    assign memory[508 ] = 16'd32520;
    assign memory[509 ] = 16'd32531;
    assign memory[510 ] = 16'd32542;
    assign memory[511 ] = 16'd32553;
    assign memory[512 ] = 16'd32564;
    assign memory[513 ] = 16'd32574;
    assign memory[514 ] = 16'd32585;
    assign memory[515 ] = 16'd32595;
    assign memory[516 ] = 16'd32605;
    assign memory[517 ] = 16'd32615;
    assign memory[518 ] = 16'd32625;
    assign memory[519 ] = 16'd32635;
    assign memory[520 ] = 16'd32644;
    assign memory[521 ] = 16'd32653;
    assign memory[522 ] = 16'd32662;
    assign memory[523 ] = 16'd32671;
    assign memory[524 ] = 16'd32679;
    assign memory[525 ] = 16'd32687;
    assign memory[526 ] = 16'd32695;
    assign memory[527 ] = 16'd32702;
    assign memory[528 ] = 16'd32709;
    assign memory[529 ] = 16'd32716;
    assign memory[530 ] = 16'd32723;
    assign memory[531 ] = 16'd32729;
    assign memory[532 ] = 16'd32734;
    assign memory[533 ] = 16'd32740;
    assign memory[534 ] = 16'd32745;
    assign memory[535 ] = 16'd32749;
    assign memory[536 ] = 16'd32753;
    assign memory[537 ] = 16'd32756;
    assign memory[538 ] = 16'd32759;
    assign memory[539 ] = 16'd32762;
    assign memory[540 ] = 16'd32764;
    assign memory[541 ] = 16'd32765;
    assign memory[542 ] = 16'd32766;
    assign memory[543 ] = 16'd32767;

endmodule
