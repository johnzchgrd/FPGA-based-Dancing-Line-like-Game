module image_reader (
    input clk,
    input valid,
    input type,
    input [1:0] song,
    input [4:0] x, y,
	output [11:0] dout
    );

    wire [12:0] ir_in;
    assign ir_in = {song, type, y, x};
    image_rom ir(clk, ir_in, dout);

endmodule

module image_rom (
    input clk,
    input [12:0] in,
    output reg [11:0] dout
    );
    
    wire [11:0] memory [8191:0];
    
    always @(posedge clk) begin
        dout = memory[in];
    end
    
    assign memory[0   ] = 12'h543;
    assign memory[1   ] = 12'h543;
    assign memory[2   ] = 12'h543;
    assign memory[3   ] = 12'h543;
    assign memory[4   ] = 12'h543;
    assign memory[5   ] = 12'h764;
    assign memory[6   ] = 12'h764;
    assign memory[7   ] = 12'h543;
    assign memory[8   ] = 12'h543;
    assign memory[9   ] = 12'h543;
    assign memory[10  ] = 12'h543;
    assign memory[11  ] = 12'h543;
    assign memory[12  ] = 12'h543;
    assign memory[13  ] = 12'h764;
    assign memory[14  ] = 12'h543;
    assign memory[15  ] = 12'h543;
    assign memory[16  ] = 12'h543;
    assign memory[17  ] = 12'h543;
    assign memory[18  ] = 12'h543;
    assign memory[19  ] = 12'h543;
    assign memory[20  ] = 12'h543;
    assign memory[21  ] = 12'h543;
    assign memory[22  ] = 12'h764;
    assign memory[23  ] = 12'h764;
    assign memory[24  ] = 12'h543;
    assign memory[25  ] = 12'h543;
    assign memory[26  ] = 12'h543;
    assign memory[27  ] = 12'h543;
    assign memory[28  ] = 12'h543;
    assign memory[29  ] = 12'h543;
    assign memory[30  ] = 12'h543;
    assign memory[31  ] = 12'h543;
    assign memory[32  ] = 12'h543;
    assign memory[33  ] = 12'h875;
    assign memory[34  ] = 12'h875;
    assign memory[35  ] = 12'h875;
    assign memory[36  ] = 12'h875;
    assign memory[37  ] = 12'h875;
    assign memory[38  ] = 12'h875;
    assign memory[39  ] = 12'h875;
    assign memory[40  ] = 12'h875;
    assign memory[41  ] = 12'h875;
    assign memory[42  ] = 12'h875;
    assign memory[43  ] = 12'h875;
    assign memory[44  ] = 12'h875;
    assign memory[45  ] = 12'ha98;
    assign memory[46  ] = 12'ha98;
    assign memory[47  ] = 12'ha98;
    assign memory[48  ] = 12'ha98;
    assign memory[49  ] = 12'ha98;
    assign memory[50  ] = 12'ha98;
    assign memory[51  ] = 12'ha98;
    assign memory[52  ] = 12'ha98;
    assign memory[53  ] = 12'h875;
    assign memory[54  ] = 12'h875;
    assign memory[55  ] = 12'h875;
    assign memory[56  ] = 12'h875;
    assign memory[57  ] = 12'h875;
    assign memory[58  ] = 12'h875;
    assign memory[59  ] = 12'h875;
    assign memory[60  ] = 12'ha98;
    assign memory[61  ] = 12'ha98;
    assign memory[62  ] = 12'ha98;
    assign memory[63  ] = 12'h543;
    assign memory[64  ] = 12'h543;
    assign memory[65  ] = 12'ha98;
    assign memory[66  ] = 12'ha98;
    assign memory[67  ] = 12'ha98;
    assign memory[68  ] = 12'ha98;
    assign memory[69  ] = 12'ha98;
    assign memory[70  ] = 12'ha98;
    assign memory[71  ] = 12'ha98;
    assign memory[72  ] = 12'ha98;
    assign memory[73  ] = 12'ha98;
    assign memory[74  ] = 12'ha98;
    assign memory[75  ] = 12'ha98;
    assign memory[76  ] = 12'ha98;
    assign memory[77  ] = 12'ha98;
    assign memory[78  ] = 12'ha98;
    assign memory[79  ] = 12'h997;
    assign memory[80  ] = 12'h997;
    assign memory[81  ] = 12'h997;
    assign memory[82  ] = 12'h997;
    assign memory[83  ] = 12'h997;
    assign memory[84  ] = 12'ha98;
    assign memory[85  ] = 12'ha98;
    assign memory[86  ] = 12'ha98;
    assign memory[87  ] = 12'ha98;
    assign memory[88  ] = 12'ha98;
    assign memory[89  ] = 12'ha98;
    assign memory[90  ] = 12'ha98;
    assign memory[91  ] = 12'ha98;
    assign memory[92  ] = 12'ha98;
    assign memory[93  ] = 12'h997;
    assign memory[94  ] = 12'h986;
    assign memory[95  ] = 12'h543;
    assign memory[96  ] = 12'h543;
    assign memory[97  ] = 12'ha98;
    assign memory[98  ] = 12'ha98;
    assign memory[99  ] = 12'ha98;
    assign memory[100 ] = 12'ha98;
    assign memory[101 ] = 12'ha98;
    assign memory[102 ] = 12'ha98;
    assign memory[103 ] = 12'ha98;
    assign memory[104 ] = 12'ha98;
    assign memory[105 ] = 12'ha98;
    assign memory[106 ] = 12'ha98;
    assign memory[107 ] = 12'h997;
    assign memory[108 ] = 12'h997;
    assign memory[109 ] = 12'h997;
    assign memory[110 ] = 12'h997;
    assign memory[111 ] = 12'h997;
    assign memory[112 ] = 12'h997;
    assign memory[113 ] = 12'h997;
    assign memory[114 ] = 12'h997;
    assign memory[115 ] = 12'h997;
    assign memory[116 ] = 12'h997;
    assign memory[117 ] = 12'h997;
    assign memory[118 ] = 12'h997;
    assign memory[119 ] = 12'h997;
    assign memory[120 ] = 12'h997;
    assign memory[121 ] = 12'h997;
    assign memory[122 ] = 12'h986;
    assign memory[123 ] = 12'h986;
    assign memory[124 ] = 12'h997;
    assign memory[125 ] = 12'h997;
    assign memory[126 ] = 12'h986;
    assign memory[127 ] = 12'h543;
    assign memory[128 ] = 12'h543;
    assign memory[129 ] = 12'ha98;
    assign memory[130 ] = 12'ha98;
    assign memory[131 ] = 12'h997;
    assign memory[132 ] = 12'h997;
    assign memory[133 ] = 12'h997;
    assign memory[134 ] = 12'h997;
    assign memory[135 ] = 12'h997;
    assign memory[136 ] = 12'h997;
    assign memory[137 ] = 12'h997;
    assign memory[138 ] = 12'h997;
    assign memory[139 ] = 12'h997;
    assign memory[140 ] = 12'h997;
    assign memory[141 ] = 12'h997;
    assign memory[142 ] = 12'h986;
    assign memory[143 ] = 12'h986;
    assign memory[144 ] = 12'h997;
    assign memory[145 ] = 12'h997;
    assign memory[146 ] = 12'h997;
    assign memory[147 ] = 12'h997;
    assign memory[148 ] = 12'h997;
    assign memory[149 ] = 12'h997;
    assign memory[150 ] = 12'h997;
    assign memory[151 ] = 12'h997;
    assign memory[152 ] = 12'h986;
    assign memory[153 ] = 12'h986;
    assign memory[154 ] = 12'h986;
    assign memory[155 ] = 12'h986;
    assign memory[156 ] = 12'h997;
    assign memory[157 ] = 12'h997;
    assign memory[158 ] = 12'h986;
    assign memory[159 ] = 12'h543;
    assign memory[160 ] = 12'h543;
    assign memory[161 ] = 12'ha98;
    assign memory[162 ] = 12'ha98;
    assign memory[163 ] = 12'h997;
    assign memory[164 ] = 12'h997;
    assign memory[165 ] = 12'h997;
    assign memory[166 ] = 12'h997;
    assign memory[167 ] = 12'h986;
    assign memory[168 ] = 12'h997;
    assign memory[169 ] = 12'h997;
    assign memory[170 ] = 12'h997;
    assign memory[171 ] = 12'h997;
    assign memory[172 ] = 12'h997;
    assign memory[173 ] = 12'h997;
    assign memory[174 ] = 12'h986;
    assign memory[175 ] = 12'h986;
    assign memory[176 ] = 12'h986;
    assign memory[177 ] = 12'h986;
    assign memory[178 ] = 12'h997;
    assign memory[179 ] = 12'h997;
    assign memory[180 ] = 12'h997;
    assign memory[181 ] = 12'h997;
    assign memory[182 ] = 12'h997;
    assign memory[183 ] = 12'h997;
    assign memory[184 ] = 12'h997;
    assign memory[185 ] = 12'h986;
    assign memory[186 ] = 12'h986;
    assign memory[187 ] = 12'h986;
    assign memory[188 ] = 12'h997;
    assign memory[189 ] = 12'h997;
    assign memory[190 ] = 12'h986;
    assign memory[191 ] = 12'h543;
    assign memory[192 ] = 12'h764;
    assign memory[193 ] = 12'h875;
    assign memory[194 ] = 12'ha98;
    assign memory[195 ] = 12'h997;
    assign memory[196 ] = 12'h997;
    assign memory[197 ] = 12'h997;
    assign memory[198 ] = 12'h986;
    assign memory[199 ] = 12'h986;
    assign memory[200 ] = 12'h986;
    assign memory[201 ] = 12'h986;
    assign memory[202 ] = 12'h986;
    assign memory[203 ] = 12'h997;
    assign memory[204 ] = 12'h997;
    assign memory[205 ] = 12'h997;
    assign memory[206 ] = 12'h997;
    assign memory[207 ] = 12'h997;
    assign memory[208 ] = 12'h997;
    assign memory[209 ] = 12'h997;
    assign memory[210 ] = 12'h997;
    assign memory[211 ] = 12'h997;
    assign memory[212 ] = 12'h997;
    assign memory[213 ] = 12'h997;
    assign memory[214 ] = 12'h997;
    assign memory[215 ] = 12'h997;
    assign memory[216 ] = 12'h997;
    assign memory[217 ] = 12'h997;
    assign memory[218 ] = 12'h986;
    assign memory[219 ] = 12'h986;
    assign memory[220 ] = 12'h997;
    assign memory[221 ] = 12'h997;
    assign memory[222 ] = 12'h986;
    assign memory[223 ] = 12'h764;
    assign memory[224 ] = 12'h764;
    assign memory[225 ] = 12'h875;
    assign memory[226 ] = 12'ha98;
    assign memory[227 ] = 12'h997;
    assign memory[228 ] = 12'h997;
    assign memory[229 ] = 12'h997;
    assign memory[230 ] = 12'h986;
    assign memory[231 ] = 12'h986;
    assign memory[232 ] = 12'h997;
    assign memory[233 ] = 12'h986;
    assign memory[234 ] = 12'h997;
    assign memory[235 ] = 12'h997;
    assign memory[236 ] = 12'h997;
    assign memory[237 ] = 12'h997;
    assign memory[238 ] = 12'h997;
    assign memory[239 ] = 12'h997;
    assign memory[240 ] = 12'h997;
    assign memory[241 ] = 12'h997;
    assign memory[242 ] = 12'h997;
    assign memory[243 ] = 12'h997;
    assign memory[244 ] = 12'h997;
    assign memory[245 ] = 12'h997;
    assign memory[246 ] = 12'h997;
    assign memory[247 ] = 12'h997;
    assign memory[248 ] = 12'h997;
    assign memory[249 ] = 12'h997;
    assign memory[250 ] = 12'h997;
    assign memory[251 ] = 12'h997;
    assign memory[252 ] = 12'h997;
    assign memory[253 ] = 12'h997;
    assign memory[254 ] = 12'h986;
    assign memory[255 ] = 12'h764;
    assign memory[256 ] = 12'h543;
    assign memory[257 ] = 12'h875;
    assign memory[258 ] = 12'ha98;
    assign memory[259 ] = 12'h997;
    assign memory[260 ] = 12'h997;
    assign memory[261 ] = 12'h997;
    assign memory[262 ] = 12'h997;
    assign memory[263 ] = 12'h997;
    assign memory[264 ] = 12'h997;
    assign memory[265 ] = 12'h997;
    assign memory[266 ] = 12'h997;
    assign memory[267 ] = 12'h997;
    assign memory[268 ] = 12'h997;
    assign memory[269 ] = 12'h997;
    assign memory[270 ] = 12'h997;
    assign memory[271 ] = 12'h997;
    assign memory[272 ] = 12'h997;
    assign memory[273 ] = 12'h997;
    assign memory[274 ] = 12'h997;
    assign memory[275 ] = 12'h997;
    assign memory[276 ] = 12'h997;
    assign memory[277 ] = 12'h997;
    assign memory[278 ] = 12'h997;
    assign memory[279 ] = 12'h997;
    assign memory[280 ] = 12'h997;
    assign memory[281 ] = 12'h997;
    assign memory[282 ] = 12'h997;
    assign memory[283 ] = 12'h997;
    assign memory[284 ] = 12'h997;
    assign memory[285 ] = 12'h997;
    assign memory[286 ] = 12'h986;
    assign memory[287 ] = 12'h543;
    assign memory[288 ] = 12'h543;
    assign memory[289 ] = 12'h875;
    assign memory[290 ] = 12'ha98;
    assign memory[291 ] = 12'h987;
    assign memory[292 ] = 12'h987;
    assign memory[293 ] = 12'h987;
    assign memory[294 ] = 12'h987;
    assign memory[295 ] = 12'h997;
    assign memory[296 ] = 12'h997;
    assign memory[297 ] = 12'h997;
    assign memory[298 ] = 12'h997;
    assign memory[299 ] = 12'h997;
    assign memory[300 ] = 12'h997;
    assign memory[301 ] = 12'h987;
    assign memory[302 ] = 12'h987;
    assign memory[303 ] = 12'h987;
    assign memory[304 ] = 12'h987;
    assign memory[305 ] = 12'h987;
    assign memory[306 ] = 12'h987;
    assign memory[307 ] = 12'h987;
    assign memory[308 ] = 12'h987;
    assign memory[309 ] = 12'h987;
    assign memory[310 ] = 12'h987;
    assign memory[311 ] = 12'h987;
    assign memory[312 ] = 12'h987;
    assign memory[313 ] = 12'h987;
    assign memory[314 ] = 12'h987;
    assign memory[315 ] = 12'h987;
    assign memory[316 ] = 12'h987;
    assign memory[317 ] = 12'h987;
    assign memory[318 ] = 12'h986;
    assign memory[319 ] = 12'h543;
    assign memory[320 ] = 12'h543;
    assign memory[321 ] = 12'h875;
    assign memory[322 ] = 12'ha98;
    assign memory[323 ] = 12'h987;
    assign memory[324 ] = 12'h987;
    assign memory[325 ] = 12'h987;
    assign memory[326 ] = 12'h987;
    assign memory[327 ] = 12'h987;
    assign memory[328 ] = 12'h987;
    assign memory[329 ] = 12'h987;
    assign memory[330 ] = 12'h987;
    assign memory[331 ] = 12'h987;
    assign memory[332 ] = 12'h987;
    assign memory[333 ] = 12'h987;
    assign memory[334 ] = 12'h987;
    assign memory[335 ] = 12'h987;
    assign memory[336 ] = 12'h987;
    assign memory[337 ] = 12'h987;
    assign memory[338 ] = 12'h987;
    assign memory[339 ] = 12'h987;
    assign memory[340 ] = 12'h987;
    assign memory[341 ] = 12'h987;
    assign memory[342 ] = 12'h987;
    assign memory[343 ] = 12'h987;
    assign memory[344 ] = 12'h987;
    assign memory[345 ] = 12'h987;
    assign memory[346 ] = 12'h987;
    assign memory[347 ] = 12'h987;
    assign memory[348 ] = 12'h987;
    assign memory[349 ] = 12'h987;
    assign memory[350 ] = 12'h986;
    assign memory[351 ] = 12'h543;
    assign memory[352 ] = 12'h543;
    assign memory[353 ] = 12'h875;
    assign memory[354 ] = 12'ha98;
    assign memory[355 ] = 12'h987;
    assign memory[356 ] = 12'h986;
    assign memory[357 ] = 12'h986;
    assign memory[358 ] = 12'h987;
    assign memory[359 ] = 12'h987;
    assign memory[360 ] = 12'h987;
    assign memory[361 ] = 12'h987;
    assign memory[362 ] = 12'h987;
    assign memory[363 ] = 12'h987;
    assign memory[364 ] = 12'h987;
    assign memory[365 ] = 12'h987;
    assign memory[366 ] = 12'h987;
    assign memory[367 ] = 12'h987;
    assign memory[368 ] = 12'h987;
    assign memory[369 ] = 12'h987;
    assign memory[370 ] = 12'h987;
    assign memory[371 ] = 12'h987;
    assign memory[372 ] = 12'h987;
    assign memory[373 ] = 12'h987;
    assign memory[374 ] = 12'h987;
    assign memory[375 ] = 12'h987;
    assign memory[376 ] = 12'h986;
    assign memory[377 ] = 12'h986;
    assign memory[378 ] = 12'h986;
    assign memory[379 ] = 12'h987;
    assign memory[380 ] = 12'h987;
    assign memory[381 ] = 12'h987;
    assign memory[382 ] = 12'h986;
    assign memory[383 ] = 12'h543;
    assign memory[384 ] = 12'h543;
    assign memory[385 ] = 12'ha98;
    assign memory[386 ] = 12'ha98;
    assign memory[387 ] = 12'h987;
    assign memory[388 ] = 12'h986;
    assign memory[389 ] = 12'h986;
    assign memory[390 ] = 12'h986;
    assign memory[391 ] = 12'h986;
    assign memory[392 ] = 12'h986;
    assign memory[393 ] = 12'h987;
    assign memory[394 ] = 12'h987;
    assign memory[395 ] = 12'h987;
    assign memory[396 ] = 12'h987;
    assign memory[397 ] = 12'h986;
    assign memory[398 ] = 12'h986;
    assign memory[399 ] = 12'h987;
    assign memory[400 ] = 12'h987;
    assign memory[401 ] = 12'h986;
    assign memory[402 ] = 12'h986;
    assign memory[403 ] = 12'h986;
    assign memory[404 ] = 12'h987;
    assign memory[405 ] = 12'h987;
    assign memory[406 ] = 12'h987;
    assign memory[407 ] = 12'h986;
    assign memory[408 ] = 12'h986;
    assign memory[409 ] = 12'h986;
    assign memory[410 ] = 12'h986;
    assign memory[411 ] = 12'h987;
    assign memory[412 ] = 12'h986;
    assign memory[413 ] = 12'h986;
    assign memory[414 ] = 12'h986;
    assign memory[415 ] = 12'h543;
    assign memory[416 ] = 12'h764;
    assign memory[417 ] = 12'ha98;
    assign memory[418 ] = 12'ha98;
    assign memory[419 ] = 12'h987;
    assign memory[420 ] = 12'h986;
    assign memory[421 ] = 12'h986;
    assign memory[422 ] = 12'h986;
    assign memory[423 ] = 12'h986;
    assign memory[424 ] = 12'h986;
    assign memory[425 ] = 12'h986;
    assign memory[426 ] = 12'h986;
    assign memory[427 ] = 12'h986;
    assign memory[428 ] = 12'h986;
    assign memory[429 ] = 12'h986;
    assign memory[430 ] = 12'h986;
    assign memory[431 ] = 12'h986;
    assign memory[432 ] = 12'h986;
    assign memory[433 ] = 12'h986;
    assign memory[434 ] = 12'h986;
    assign memory[435 ] = 12'h986;
    assign memory[436 ] = 12'h986;
    assign memory[437 ] = 12'h986;
    assign memory[438 ] = 12'h987;
    assign memory[439 ] = 12'h986;
    assign memory[440 ] = 12'h986;
    assign memory[441 ] = 12'h986;
    assign memory[442 ] = 12'h986;
    assign memory[443 ] = 12'h986;
    assign memory[444 ] = 12'h986;
    assign memory[445 ] = 12'h986;
    assign memory[446 ] = 12'h986;
    assign memory[447 ] = 12'h764;
    assign memory[448 ] = 12'h543;
    assign memory[449 ] = 12'ha98;
    assign memory[450 ] = 12'ha98;
    assign memory[451 ] = 12'h986;
    assign memory[452 ] = 12'h986;
    assign memory[453 ] = 12'h986;
    assign memory[454 ] = 12'h986;
    assign memory[455 ] = 12'h986;
    assign memory[456 ] = 12'h986;
    assign memory[457 ] = 12'h986;
    assign memory[458 ] = 12'h986;
    assign memory[459 ] = 12'h986;
    assign memory[460 ] = 12'h986;
    assign memory[461 ] = 12'h986;
    assign memory[462 ] = 12'h986;
    assign memory[463 ] = 12'h986;
    assign memory[464 ] = 12'h986;
    assign memory[465 ] = 12'h986;
    assign memory[466 ] = 12'h986;
    assign memory[467 ] = 12'h986;
    assign memory[468 ] = 12'h986;
    assign memory[469 ] = 12'h986;
    assign memory[470 ] = 12'h986;
    assign memory[471 ] = 12'h986;
    assign memory[472 ] = 12'h986;
    assign memory[473 ] = 12'h986;
    assign memory[474 ] = 12'h986;
    assign memory[475 ] = 12'h986;
    assign memory[476 ] = 12'h543;
    assign memory[477 ] = 12'h543;
    assign memory[478 ] = 12'h543;
    assign memory[479 ] = 12'h543;
    assign memory[480 ] = 12'h543;
    assign memory[481 ] = 12'h543;
    assign memory[482 ] = 12'h543;
    assign memory[483 ] = 12'h543;
    assign memory[484 ] = 12'h543;
    assign memory[485 ] = 12'h543;
    assign memory[486 ] = 12'h543;
    assign memory[487 ] = 12'h543;
    assign memory[488 ] = 12'h543;
    assign memory[489 ] = 12'h543;
    assign memory[490 ] = 12'h764;
    assign memory[491 ] = 12'h543;
    assign memory[492 ] = 12'h543;
    assign memory[493 ] = 12'h543;
    assign memory[494 ] = 12'h543;
    assign memory[495 ] = 12'h543;
    assign memory[496 ] = 12'h543;
    assign memory[497 ] = 12'h543;
    assign memory[498 ] = 12'h543;
    assign memory[499 ] = 12'h543;
    assign memory[500 ] = 12'h543;
    assign memory[501 ] = 12'h543;
    assign memory[502 ] = 12'h543;
    assign memory[503 ] = 12'h543;
    assign memory[504 ] = 12'h543;
    assign memory[505 ] = 12'h764;
    assign memory[506 ] = 12'h764;
    assign memory[507 ] = 12'h543;
    assign memory[508 ] = 12'h543;
    assign memory[509 ] = 12'h543;
    assign memory[510 ] = 12'h543;
    assign memory[511 ] = 12'h543;
    assign memory[512 ] = 12'h543;
    assign memory[513 ] = 12'h543;
    assign memory[514 ] = 12'h543;
    assign memory[515 ] = 12'h543;
    assign memory[516 ] = 12'h543;
    assign memory[517 ] = 12'h543;
    assign memory[518 ] = 12'h543;
    assign memory[519 ] = 12'h543;
    assign memory[520 ] = 12'h543;
    assign memory[521 ] = 12'h543;
    assign memory[522 ] = 12'h764;
    assign memory[523 ] = 12'h543;
    assign memory[524 ] = 12'h543;
    assign memory[525 ] = 12'h543;
    assign memory[526 ] = 12'h543;
    assign memory[527 ] = 12'h543;
    assign memory[528 ] = 12'h543;
    assign memory[529 ] = 12'h543;
    assign memory[530 ] = 12'h543;
    assign memory[531 ] = 12'h543;
    assign memory[532 ] = 12'h543;
    assign memory[533 ] = 12'h543;
    assign memory[534 ] = 12'h543;
    assign memory[535 ] = 12'h543;
    assign memory[536 ] = 12'h543;
    assign memory[537 ] = 12'h764;
    assign memory[538 ] = 12'h764;
    assign memory[539 ] = 12'h543;
    assign memory[540 ] = 12'h543;
    assign memory[541 ] = 12'h543;
    assign memory[542 ] = 12'h543;
    assign memory[543 ] = 12'h543;
    assign memory[544 ] = 12'ha98;
    assign memory[545 ] = 12'ha98;
    assign memory[546 ] = 12'ha98;
    assign memory[547 ] = 12'ha98;
    assign memory[548 ] = 12'ha98;
    assign memory[549 ] = 12'ha98;
    assign memory[550 ] = 12'ha98;
    assign memory[551 ] = 12'ha98;
    assign memory[552 ] = 12'ha98;
    assign memory[553 ] = 12'ha98;
    assign memory[554 ] = 12'ha98;
    assign memory[555 ] = 12'ha98;
    assign memory[556 ] = 12'ha98;
    assign memory[557 ] = 12'ha98;
    assign memory[558 ] = 12'h875;
    assign memory[559 ] = 12'h543;
    assign memory[560 ] = 12'h543;
    assign memory[561 ] = 12'h875;
    assign memory[562 ] = 12'h875;
    assign memory[563 ] = 12'ha98;
    assign memory[564 ] = 12'ha98;
    assign memory[565 ] = 12'ha98;
    assign memory[566 ] = 12'ha98;
    assign memory[567 ] = 12'ha98;
    assign memory[568 ] = 12'ha98;
    assign memory[569 ] = 12'ha98;
    assign memory[570 ] = 12'ha98;
    assign memory[571 ] = 12'ha98;
    assign memory[572 ] = 12'ha98;
    assign memory[573 ] = 12'ha98;
    assign memory[574 ] = 12'ha98;
    assign memory[575 ] = 12'ha98;
    assign memory[576 ] = 12'ha98;
    assign memory[577 ] = 12'h997;
    assign memory[578 ] = 12'h997;
    assign memory[579 ] = 12'h997;
    assign memory[580 ] = 12'h997;
    assign memory[581 ] = 12'h997;
    assign memory[582 ] = 12'h997;
    assign memory[583 ] = 12'h997;
    assign memory[584 ] = 12'h997;
    assign memory[585 ] = 12'h997;
    assign memory[586 ] = 12'h997;
    assign memory[587 ] = 12'h997;
    assign memory[588 ] = 12'h997;
    assign memory[589 ] = 12'h997;
    assign memory[590 ] = 12'h986;
    assign memory[591 ] = 12'h543;
    assign memory[592 ] = 12'h543;
    assign memory[593 ] = 12'ha98;
    assign memory[594 ] = 12'ha98;
    assign memory[595 ] = 12'ha98;
    assign memory[596 ] = 12'ha98;
    assign memory[597 ] = 12'ha98;
    assign memory[598 ] = 12'ha98;
    assign memory[599 ] = 12'ha98;
    assign memory[600 ] = 12'ha98;
    assign memory[601 ] = 12'ha98;
    assign memory[602 ] = 12'ha98;
    assign memory[603 ] = 12'ha98;
    assign memory[604 ] = 12'ha98;
    assign memory[605 ] = 12'ha98;
    assign memory[606 ] = 12'ha98;
    assign memory[607 ] = 12'ha98;
    assign memory[608 ] = 12'h997;
    assign memory[609 ] = 12'h997;
    assign memory[610 ] = 12'h997;
    assign memory[611 ] = 12'h997;
    assign memory[612 ] = 12'h997;
    assign memory[613 ] = 12'h997;
    assign memory[614 ] = 12'h997;
    assign memory[615 ] = 12'h997;
    assign memory[616 ] = 12'h997;
    assign memory[617 ] = 12'h986;
    assign memory[618 ] = 12'h997;
    assign memory[619 ] = 12'h997;
    assign memory[620 ] = 12'h997;
    assign memory[621 ] = 12'h997;
    assign memory[622 ] = 12'h986;
    assign memory[623 ] = 12'h543;
    assign memory[624 ] = 12'h543;
    assign memory[625 ] = 12'ha98;
    assign memory[626 ] = 12'ha98;
    assign memory[627 ] = 12'h997;
    assign memory[628 ] = 12'h997;
    assign memory[629 ] = 12'h997;
    assign memory[630 ] = 12'h997;
    assign memory[631 ] = 12'h997;
    assign memory[632 ] = 12'h997;
    assign memory[633 ] = 12'h997;
    assign memory[634 ] = 12'h997;
    assign memory[635 ] = 12'h997;
    assign memory[636 ] = 12'h997;
    assign memory[637 ] = 12'h997;
    assign memory[638 ] = 12'h997;
    assign memory[639 ] = 12'h997;
    assign memory[640 ] = 12'h997;
    assign memory[641 ] = 12'h997;
    assign memory[642 ] = 12'h997;
    assign memory[643 ] = 12'h997;
    assign memory[644 ] = 12'h997;
    assign memory[645 ] = 12'h997;
    assign memory[646 ] = 12'h986;
    assign memory[647 ] = 12'h986;
    assign memory[648 ] = 12'h986;
    assign memory[649 ] = 12'h986;
    assign memory[650 ] = 12'h986;
    assign memory[651 ] = 12'h997;
    assign memory[652 ] = 12'h997;
    assign memory[653 ] = 12'h997;
    assign memory[654 ] = 12'h986;
    assign memory[655 ] = 12'h764;
    assign memory[656 ] = 12'h764;
    assign memory[657 ] = 12'ha98;
    assign memory[658 ] = 12'ha98;
    assign memory[659 ] = 12'h997;
    assign memory[660 ] = 12'h997;
    assign memory[661 ] = 12'h997;
    assign memory[662 ] = 12'h997;
    assign memory[663 ] = 12'h997;
    assign memory[664 ] = 12'h997;
    assign memory[665 ] = 12'h986;
    assign memory[666 ] = 12'h997;
    assign memory[667 ] = 12'h997;
    assign memory[668 ] = 12'h997;
    assign memory[669 ] = 12'h997;
    assign memory[670 ] = 12'h997;
    assign memory[671 ] = 12'h997;
    assign memory[672 ] = 12'h986;
    assign memory[673 ] = 12'h986;
    assign memory[674 ] = 12'h997;
    assign memory[675 ] = 12'h997;
    assign memory[676 ] = 12'h997;
    assign memory[677 ] = 12'h997;
    assign memory[678 ] = 12'h997;
    assign memory[679 ] = 12'h997;
    assign memory[680 ] = 12'h986;
    assign memory[681 ] = 12'h986;
    assign memory[682 ] = 12'h986;
    assign memory[683 ] = 12'h997;
    assign memory[684 ] = 12'h997;
    assign memory[685 ] = 12'h997;
    assign memory[686 ] = 12'h986;
    assign memory[687 ] = 12'h764;
    assign memory[688 ] = 12'h764;
    assign memory[689 ] = 12'ha98;
    assign memory[690 ] = 12'ha98;
    assign memory[691 ] = 12'h997;
    assign memory[692 ] = 12'h986;
    assign memory[693 ] = 12'h986;
    assign memory[694 ] = 12'h997;
    assign memory[695 ] = 12'h997;
    assign memory[696 ] = 12'h997;
    assign memory[697 ] = 12'h997;
    assign memory[698 ] = 12'h997;
    assign memory[699 ] = 12'h997;
    assign memory[700 ] = 12'h997;
    assign memory[701 ] = 12'h986;
    assign memory[702 ] = 12'h986;
    assign memory[703 ] = 12'h986;
    assign memory[704 ] = 12'h986;
    assign memory[705 ] = 12'h986;
    assign memory[706 ] = 12'h997;
    assign memory[707 ] = 12'h997;
    assign memory[708 ] = 12'h997;
    assign memory[709 ] = 12'h997;
    assign memory[710 ] = 12'h997;
    assign memory[711 ] = 12'h997;
    assign memory[712 ] = 12'h997;
    assign memory[713 ] = 12'h997;
    assign memory[714 ] = 12'h997;
    assign memory[715 ] = 12'h997;
    assign memory[716 ] = 12'h997;
    assign memory[717 ] = 12'h997;
    assign memory[718 ] = 12'h986;
    assign memory[719 ] = 12'h543;
    assign memory[720 ] = 12'h543;
    assign memory[721 ] = 12'ha98;
    assign memory[722 ] = 12'ha98;
    assign memory[723 ] = 12'h997;
    assign memory[724 ] = 12'h986;
    assign memory[725 ] = 12'h986;
    assign memory[726 ] = 12'h986;
    assign memory[727 ] = 12'h997;
    assign memory[728 ] = 12'h997;
    assign memory[729 ] = 12'h997;
    assign memory[730 ] = 12'h997;
    assign memory[731 ] = 12'h997;
    assign memory[732 ] = 12'h997;
    assign memory[733 ] = 12'h997;
    assign memory[734 ] = 12'h986;
    assign memory[735 ] = 12'h986;
    assign memory[736 ] = 12'h997;
    assign memory[737 ] = 12'h997;
    assign memory[738 ] = 12'h997;
    assign memory[739 ] = 12'h997;
    assign memory[740 ] = 12'h997;
    assign memory[741 ] = 12'h997;
    assign memory[742 ] = 12'h997;
    assign memory[743 ] = 12'h997;
    assign memory[744 ] = 12'h997;
    assign memory[745 ] = 12'h997;
    assign memory[746 ] = 12'h997;
    assign memory[747 ] = 12'h997;
    assign memory[748 ] = 12'h997;
    assign memory[749 ] = 12'h997;
    assign memory[750 ] = 12'h986;
    assign memory[751 ] = 12'h543;
    assign memory[752 ] = 12'h543;
    assign memory[753 ] = 12'ha98;
    assign memory[754 ] = 12'ha98;
    assign memory[755 ] = 12'h997;
    assign memory[756 ] = 12'h997;
    assign memory[757 ] = 12'h986;
    assign memory[758 ] = 12'h997;
    assign memory[759 ] = 12'h997;
    assign memory[760 ] = 12'h997;
    assign memory[761 ] = 12'h997;
    assign memory[762 ] = 12'h997;
    assign memory[763 ] = 12'h997;
    assign memory[764 ] = 12'h997;
    assign memory[765 ] = 12'h997;
    assign memory[766 ] = 12'h997;
    assign memory[767 ] = 12'h997;
    assign memory[768 ] = 12'h997;
    assign memory[769 ] = 12'h997;
    assign memory[770 ] = 12'h987;
    assign memory[771 ] = 12'h987;
    assign memory[772 ] = 12'h987;
    assign memory[773 ] = 12'h987;
    assign memory[774 ] = 12'h987;
    assign memory[775 ] = 12'h987;
    assign memory[776 ] = 12'h987;
    assign memory[777 ] = 12'h987;
    assign memory[778 ] = 12'h997;
    assign memory[779 ] = 12'h997;
    assign memory[780 ] = 12'h997;
    assign memory[781 ] = 12'h997;
    assign memory[782 ] = 12'h986;
    assign memory[783 ] = 12'h543;
    assign memory[784 ] = 12'h543;
    assign memory[785 ] = 12'ha98;
    assign memory[786 ] = 12'ha98;
    assign memory[787 ] = 12'h997;
    assign memory[788 ] = 12'h997;
    assign memory[789 ] = 12'h997;
    assign memory[790 ] = 12'h997;
    assign memory[791 ] = 12'h997;
    assign memory[792 ] = 12'h997;
    assign memory[793 ] = 12'h997;
    assign memory[794 ] = 12'h997;
    assign memory[795 ] = 12'h997;
    assign memory[796 ] = 12'h997;
    assign memory[797 ] = 12'h997;
    assign memory[798 ] = 12'h997;
    assign memory[799 ] = 12'h997;
    assign memory[800 ] = 12'h987;
    assign memory[801 ] = 12'h987;
    assign memory[802 ] = 12'h987;
    assign memory[803 ] = 12'h987;
    assign memory[804 ] = 12'h987;
    assign memory[805 ] = 12'h987;
    assign memory[806 ] = 12'h987;
    assign memory[807 ] = 12'h987;
    assign memory[808 ] = 12'h987;
    assign memory[809 ] = 12'h987;
    assign memory[810 ] = 12'h987;
    assign memory[811 ] = 12'h987;
    assign memory[812 ] = 12'h987;
    assign memory[813 ] = 12'h987;
    assign memory[814 ] = 12'h986;
    assign memory[815 ] = 12'h543;
    assign memory[816 ] = 12'h543;
    assign memory[817 ] = 12'ha98;
    assign memory[818 ] = 12'ha98;
    assign memory[819 ] = 12'h997;
    assign memory[820 ] = 12'h987;
    assign memory[821 ] = 12'h987;
    assign memory[822 ] = 12'h987;
    assign memory[823 ] = 12'h987;
    assign memory[824 ] = 12'h987;
    assign memory[825 ] = 12'h987;
    assign memory[826 ] = 12'h987;
    assign memory[827 ] = 12'h997;
    assign memory[828 ] = 12'h997;
    assign memory[829 ] = 12'h997;
    assign memory[830 ] = 12'h997;
    assign memory[831 ] = 12'h987;
    assign memory[832 ] = 12'h987;
    assign memory[833 ] = 12'h987;
    assign memory[834 ] = 12'h987;
    assign memory[835 ] = 12'h986;
    assign memory[836 ] = 12'h986;
    assign memory[837 ] = 12'h987;
    assign memory[838 ] = 12'h987;
    assign memory[839 ] = 12'h987;
    assign memory[840 ] = 12'h987;
    assign memory[841 ] = 12'h987;
    assign memory[842 ] = 12'h987;
    assign memory[843 ] = 12'h987;
    assign memory[844 ] = 12'h987;
    assign memory[845 ] = 12'h987;
    assign memory[846 ] = 12'h986;
    assign memory[847 ] = 12'h543;
    assign memory[848 ] = 12'h543;
    assign memory[849 ] = 12'ha98;
    assign memory[850 ] = 12'ha98;
    assign memory[851 ] = 12'h987;
    assign memory[852 ] = 12'h987;
    assign memory[853 ] = 12'h987;
    assign memory[854 ] = 12'h987;
    assign memory[855 ] = 12'h987;
    assign memory[856 ] = 12'h987;
    assign memory[857 ] = 12'h987;
    assign memory[858 ] = 12'h987;
    assign memory[859 ] = 12'h986;
    assign memory[860 ] = 12'h986;
    assign memory[861 ] = 12'h987;
    assign memory[862 ] = 12'h987;
    assign memory[863 ] = 12'h987;
    assign memory[864 ] = 12'h987;
    assign memory[865 ] = 12'h986;
    assign memory[866 ] = 12'h986;
    assign memory[867 ] = 12'h986;
    assign memory[868 ] = 12'h986;
    assign memory[869 ] = 12'h986;
    assign memory[870 ] = 12'h987;
    assign memory[871 ] = 12'h987;
    assign memory[872 ] = 12'h987;
    assign memory[873 ] = 12'h987;
    assign memory[874 ] = 12'h987;
    assign memory[875 ] = 12'h987;
    assign memory[876 ] = 12'h987;
    assign memory[877 ] = 12'h987;
    assign memory[878 ] = 12'h986;
    assign memory[879 ] = 12'h764;
    assign memory[880 ] = 12'h764;
    assign memory[881 ] = 12'ha98;
    assign memory[882 ] = 12'ha98;
    assign memory[883 ] = 12'h987;
    assign memory[884 ] = 12'h987;
    assign memory[885 ] = 12'h987;
    assign memory[886 ] = 12'h987;
    assign memory[887 ] = 12'h987;
    assign memory[888 ] = 12'h987;
    assign memory[889 ] = 12'h986;
    assign memory[890 ] = 12'h986;
    assign memory[891 ] = 12'h986;
    assign memory[892 ] = 12'h986;
    assign memory[893 ] = 12'h986;
    assign memory[894 ] = 12'h987;
    assign memory[895 ] = 12'h987;
    assign memory[896 ] = 12'h986;
    assign memory[897 ] = 12'h986;
    assign memory[898 ] = 12'h986;
    assign memory[899 ] = 12'h986;
    assign memory[900 ] = 12'h986;
    assign memory[901 ] = 12'h986;
    assign memory[902 ] = 12'h987;
    assign memory[903 ] = 12'h987;
    assign memory[904 ] = 12'h987;
    assign memory[905 ] = 12'h987;
    assign memory[906 ] = 12'h987;
    assign memory[907 ] = 12'h986;
    assign memory[908 ] = 12'h986;
    assign memory[909 ] = 12'h986;
    assign memory[910 ] = 12'h986;
    assign memory[911 ] = 12'h543;
    assign memory[912 ] = 12'h543;
    assign memory[913 ] = 12'ha98;
    assign memory[914 ] = 12'ha98;
    assign memory[915 ] = 12'h987;
    assign memory[916 ] = 12'h987;
    assign memory[917 ] = 12'h987;
    assign memory[918 ] = 12'h987;
    assign memory[919 ] = 12'h987;
    assign memory[920 ] = 12'h986;
    assign memory[921 ] = 12'h986;
    assign memory[922 ] = 12'h986;
    assign memory[923 ] = 12'h986;
    assign memory[924 ] = 12'h986;
    assign memory[925 ] = 12'h986;
    assign memory[926 ] = 12'h986;
    assign memory[927 ] = 12'h986;
    assign memory[928 ] = 12'h986;
    assign memory[929 ] = 12'h986;
    assign memory[930 ] = 12'h986;
    assign memory[931 ] = 12'h986;
    assign memory[932 ] = 12'h986;
    assign memory[933 ] = 12'h986;
    assign memory[934 ] = 12'h987;
    assign memory[935 ] = 12'h987;
    assign memory[936 ] = 12'h986;
    assign memory[937 ] = 12'h986;
    assign memory[938 ] = 12'h986;
    assign memory[939 ] = 12'h986;
    assign memory[940 ] = 12'h986;
    assign memory[941 ] = 12'h986;
    assign memory[942 ] = 12'h875;
    assign memory[943 ] = 12'h543;
    assign memory[944 ] = 12'h543;
    assign memory[945 ] = 12'h543;
    assign memory[946 ] = 12'ha98;
    assign memory[947 ] = 12'h987;
    assign memory[948 ] = 12'h987;
    assign memory[949 ] = 12'h987;
    assign memory[950 ] = 12'h986;
    assign memory[951 ] = 12'h986;
    assign memory[952 ] = 12'h986;
    assign memory[953 ] = 12'h986;
    assign memory[954 ] = 12'h986;
    assign memory[955 ] = 12'h986;
    assign memory[956 ] = 12'h986;
    assign memory[957 ] = 12'h986;
    assign memory[958 ] = 12'h986;
    assign memory[959 ] = 12'h986;
    assign memory[960 ] = 12'h875;
    assign memory[961 ] = 12'h875;
    assign memory[962 ] = 12'h875;
    assign memory[963 ] = 12'h875;
    assign memory[964 ] = 12'h875;
    assign memory[965 ] = 12'h986;
    assign memory[966 ] = 12'h986;
    assign memory[967 ] = 12'h986;
    assign memory[968 ] = 12'h986;
    assign memory[969 ] = 12'h986;
    assign memory[970 ] = 12'h986;
    assign memory[971 ] = 12'h986;
    assign memory[972 ] = 12'h986;
    assign memory[973 ] = 12'h986;
    assign memory[974 ] = 12'h875;
    assign memory[975 ] = 12'h543;
    assign memory[976 ] = 12'h543;
    assign memory[977 ] = 12'h543;
    assign memory[978 ] = 12'ha98;
    assign memory[979 ] = 12'h986;
    assign memory[980 ] = 12'h986;
    assign memory[981 ] = 12'h986;
    assign memory[982 ] = 12'h986;
    assign memory[983 ] = 12'h986;
    assign memory[984 ] = 12'h875;
    assign memory[985 ] = 12'h875;
    assign memory[986 ] = 12'h875;
    assign memory[987 ] = 12'h875;
    assign memory[988 ] = 12'h875;
    assign memory[989 ] = 12'h875;
    assign memory[990 ] = 12'h875;
    assign memory[991 ] = 12'h986;
    assign memory[992 ] = 12'h543;
    assign memory[993 ] = 12'h543;
    assign memory[994 ] = 12'h543;
    assign memory[995 ] = 12'h543;
    assign memory[996 ] = 12'h543;
    assign memory[997 ] = 12'h764;
    assign memory[998 ] = 12'h764;
    assign memory[999 ] = 12'h543;
    assign memory[1000] = 12'h543;
    assign memory[1001] = 12'h543;
    assign memory[1002] = 12'h543;
    assign memory[1003] = 12'h543;
    assign memory[1004] = 12'h543;
    assign memory[1005] = 12'h764;
    assign memory[1006] = 12'h543;
    assign memory[1007] = 12'h543;
    assign memory[1008] = 12'h543;
    assign memory[1009] = 12'h543;
    assign memory[1010] = 12'h543;
    assign memory[1011] = 12'h543;
    assign memory[1012] = 12'h543;
    assign memory[1013] = 12'h543;
    assign memory[1014] = 12'h764;
    assign memory[1015] = 12'h764;
    assign memory[1016] = 12'h543;
    assign memory[1017] = 12'h543;
    assign memory[1018] = 12'h543;
    assign memory[1019] = 12'h543;
    assign memory[1020] = 12'h543;
    assign memory[1021] = 12'h543;
    assign memory[1022] = 12'h543;
    assign memory[1023] = 12'h543;
    assign memory[1024] = 12'h998;
    assign memory[1025] = 12'h898;
    assign memory[1026] = 12'h888;
    assign memory[1027] = 12'h998;
    assign memory[1028] = 12'h888;
    assign memory[1029] = 12'h888;
    assign memory[1030] = 12'h888;
    assign memory[1031] = 12'h887;
    assign memory[1032] = 12'h887;
    assign memory[1033] = 12'h998;
    assign memory[1034] = 12'h888;
    assign memory[1035] = 12'h998;
    assign memory[1036] = 12'h998;
    assign memory[1037] = 12'h888;
    assign memory[1038] = 12'h898;
    assign memory[1039] = 12'h888;
    assign memory[1040] = 12'h998;
    assign memory[1041] = 12'h998;
    assign memory[1042] = 12'h999;
    assign memory[1043] = 12'h998;
    assign memory[1044] = 12'h998;
    assign memory[1045] = 12'h999;
    assign memory[1046] = 12'h998;
    assign memory[1047] = 12'h888;
    assign memory[1048] = 12'h888;
    assign memory[1049] = 12'h998;
    assign memory[1050] = 12'h998;
    assign memory[1051] = 12'h887;
    assign memory[1052] = 12'h998;
    assign memory[1053] = 12'h998;
    assign memory[1054] = 12'h888;
    assign memory[1055] = 12'h998;
    assign memory[1056] = 12'h888;
    assign memory[1057] = 12'h998;
    assign memory[1058] = 12'h998;
    assign memory[1059] = 12'h888;
    assign memory[1060] = 12'h998;
    assign memory[1061] = 12'h887;
    assign memory[1062] = 12'h998;
    assign memory[1063] = 12'h998;
    assign memory[1064] = 12'h998;
    assign memory[1065] = 12'h888;
    assign memory[1066] = 12'h888;
    assign memory[1067] = 12'h998;
    assign memory[1068] = 12'h999;
    assign memory[1069] = 12'h998;
    assign memory[1070] = 12'h998;
    assign memory[1071] = 12'h888;
    assign memory[1072] = 12'h999;
    assign memory[1073] = 12'h998;
    assign memory[1074] = 12'h999;
    assign memory[1075] = 12'h999;
    assign memory[1076] = 12'h998;
    assign memory[1077] = 12'h998;
    assign memory[1078] = 12'h998;
    assign memory[1079] = 12'h999;
    assign memory[1080] = 12'h998;
    assign memory[1081] = 12'h998;
    assign memory[1082] = 12'h998;
    assign memory[1083] = 12'h998;
    assign memory[1084] = 12'h999;
    assign memory[1085] = 12'h998;
    assign memory[1086] = 12'h999;
    assign memory[1087] = 12'h898;
    assign memory[1088] = 12'h888;
    assign memory[1089] = 12'h888;
    assign memory[1090] = 12'h998;
    assign memory[1091] = 12'h888;
    assign memory[1092] = 12'h998;
    assign memory[1093] = 12'h888;
    assign memory[1094] = 12'h998;
    assign memory[1095] = 12'h998;
    assign memory[1096] = 12'h998;
    assign memory[1097] = 12'h998;
    assign memory[1098] = 12'h888;
    assign memory[1099] = 12'h998;
    assign memory[1100] = 12'h888;
    assign memory[1101] = 12'h887;
    assign memory[1102] = 12'h888;
    assign memory[1103] = 12'h999;
    assign memory[1104] = 12'h998;
    assign memory[1105] = 12'h998;
    assign memory[1106] = 12'h998;
    assign memory[1107] = 12'h998;
    assign memory[1108] = 12'h888;
    assign memory[1109] = 12'h999;
    assign memory[1110] = 12'h998;
    assign memory[1111] = 12'h998;
    assign memory[1112] = 12'h998;
    assign memory[1113] = 12'h999;
    assign memory[1114] = 12'h998;
    assign memory[1115] = 12'h898;
    assign memory[1116] = 12'h998;
    assign memory[1117] = 12'h888;
    assign memory[1118] = 12'h998;
    assign memory[1119] = 12'h998;
    assign memory[1120] = 12'h888;
    assign memory[1121] = 12'h887;
    assign memory[1122] = 12'h998;
    assign memory[1123] = 12'h998;
    assign memory[1124] = 12'h998;
    assign memory[1125] = 12'h888;
    assign memory[1126] = 12'h898;
    assign memory[1127] = 12'h999;
    assign memory[1128] = 12'h998;
    assign memory[1129] = 12'h998;
    assign memory[1130] = 12'h998;
    assign memory[1131] = 12'h888;
    assign memory[1132] = 12'h998;
    assign memory[1133] = 12'h998;
    assign memory[1134] = 12'h999;
    assign memory[1135] = 12'h998;
    assign memory[1136] = 12'h998;
    assign memory[1137] = 12'h999;
    assign memory[1138] = 12'h888;
    assign memory[1139] = 12'h888;
    assign memory[1140] = 12'h998;
    assign memory[1141] = 12'h888;
    assign memory[1142] = 12'h998;
    assign memory[1143] = 12'h998;
    assign memory[1144] = 12'h998;
    assign memory[1145] = 12'h998;
    assign memory[1146] = 12'h998;
    assign memory[1147] = 12'h888;
    assign memory[1148] = 12'h888;
    assign memory[1149] = 12'h999;
    assign memory[1150] = 12'h999;
    assign memory[1151] = 12'h998;
    assign memory[1152] = 12'h998;
    assign memory[1153] = 12'h998;
    assign memory[1154] = 12'h998;
    assign memory[1155] = 12'h998;
    assign memory[1156] = 12'h998;
    assign memory[1157] = 12'h898;
    assign memory[1158] = 12'h898;
    assign memory[1159] = 12'h998;
    assign memory[1160] = 12'h888;
    assign memory[1161] = 12'h998;
    assign memory[1162] = 12'h998;
    assign memory[1163] = 12'h998;
    assign memory[1164] = 12'h998;
    assign memory[1165] = 12'h998;
    assign memory[1166] = 12'h999;
    assign memory[1167] = 12'h998;
    assign memory[1168] = 12'h998;
    assign memory[1169] = 12'h998;
    assign memory[1170] = 12'h998;
    assign memory[1171] = 12'h999;
    assign memory[1172] = 12'h888;
    assign memory[1173] = 12'h998;
    assign memory[1174] = 12'h887;
    assign memory[1175] = 12'h888;
    assign memory[1176] = 12'h998;
    assign memory[1177] = 12'h998;
    assign memory[1178] = 12'h998;
    assign memory[1179] = 12'h898;
    assign memory[1180] = 12'h998;
    assign memory[1181] = 12'h998;
    assign memory[1182] = 12'h998;
    assign memory[1183] = 12'h998;
    assign memory[1184] = 12'h998;
    assign memory[1185] = 12'h888;
    assign memory[1186] = 12'h998;
    assign memory[1187] = 12'h888;
    assign memory[1188] = 12'h998;
    assign memory[1189] = 12'h998;
    assign memory[1190] = 12'h998;
    assign memory[1191] = 12'h998;
    assign memory[1192] = 12'h898;
    assign memory[1193] = 12'h888;
    assign memory[1194] = 12'h999;
    assign memory[1195] = 12'h998;
    assign memory[1196] = 12'h888;
    assign memory[1197] = 12'h888;
    assign memory[1198] = 12'h998;
    assign memory[1199] = 12'h998;
    assign memory[1200] = 12'h999;
    assign memory[1201] = 12'h998;
    assign memory[1202] = 12'h998;
    assign memory[1203] = 12'h998;
    assign memory[1204] = 12'h887;
    assign memory[1205] = 12'h998;
    assign memory[1206] = 12'h998;
    assign memory[1207] = 12'h998;
    assign memory[1208] = 12'h888;
    assign memory[1209] = 12'h888;
    assign memory[1210] = 12'h998;
    assign memory[1211] = 12'h998;
    assign memory[1212] = 12'h998;
    assign memory[1213] = 12'h888;
    assign memory[1214] = 12'h888;
    assign memory[1215] = 12'h999;
    assign memory[1216] = 12'h998;
    assign memory[1217] = 12'h999;
    assign memory[1218] = 12'h888;
    assign memory[1219] = 12'h998;
    assign memory[1220] = 12'h998;
    assign memory[1221] = 12'h998;
    assign memory[1222] = 12'h998;
    assign memory[1223] = 12'h898;
    assign memory[1224] = 12'h888;
    assign memory[1225] = 12'h999;
    assign memory[1226] = 12'h888;
    assign memory[1227] = 12'h888;
    assign memory[1228] = 12'h999;
    assign memory[1229] = 12'h888;
    assign memory[1230] = 12'h898;
    assign memory[1231] = 12'h998;
    assign memory[1232] = 12'h999;
    assign memory[1233] = 12'h887;
    assign memory[1234] = 12'h998;
    assign memory[1235] = 12'h998;
    assign memory[1236] = 12'h888;
    assign memory[1237] = 12'h998;
    assign memory[1238] = 12'h888;
    assign memory[1239] = 12'h998;
    assign memory[1240] = 12'h888;
    assign memory[1241] = 12'h998;
    assign memory[1242] = 12'h888;
    assign memory[1243] = 12'h998;
    assign memory[1244] = 12'h999;
    assign memory[1245] = 12'h998;
    assign memory[1246] = 12'h998;
    assign memory[1247] = 12'h998;
    assign memory[1248] = 12'h888;
    assign memory[1249] = 12'h998;
    assign memory[1250] = 12'h998;
    assign memory[1251] = 12'h888;
    assign memory[1252] = 12'h998;
    assign memory[1253] = 12'h998;
    assign memory[1254] = 12'h998;
    assign memory[1255] = 12'h998;
    assign memory[1256] = 12'h998;
    assign memory[1257] = 12'h999;
    assign memory[1258] = 12'h888;
    assign memory[1259] = 12'h998;
    assign memory[1260] = 12'h999;
    assign memory[1261] = 12'h998;
    assign memory[1262] = 12'h998;
    assign memory[1263] = 12'h888;
    assign memory[1264] = 12'h998;
    assign memory[1265] = 12'h999;
    assign memory[1266] = 12'h999;
    assign memory[1267] = 12'h888;
    assign memory[1268] = 12'h999;
    assign memory[1269] = 12'h887;
    assign memory[1270] = 12'h999;
    assign memory[1271] = 12'h999;
    assign memory[1272] = 12'h888;
    assign memory[1273] = 12'h998;
    assign memory[1274] = 12'h999;
    assign memory[1275] = 12'h998;
    assign memory[1276] = 12'h998;
    assign memory[1277] = 12'h998;
    assign memory[1278] = 12'h998;
    assign memory[1279] = 12'h998;
    assign memory[1280] = 12'h998;
    assign memory[1281] = 12'h888;
    assign memory[1282] = 12'h998;
    assign memory[1283] = 12'h888;
    assign memory[1284] = 12'h999;
    assign memory[1285] = 12'h888;
    assign memory[1286] = 12'h888;
    assign memory[1287] = 12'h998;
    assign memory[1288] = 12'h888;
    assign memory[1289] = 12'h888;
    assign memory[1290] = 12'h887;
    assign memory[1291] = 12'h888;
    assign memory[1292] = 12'h998;
    assign memory[1293] = 12'h998;
    assign memory[1294] = 12'h888;
    assign memory[1295] = 12'h999;
    assign memory[1296] = 12'h999;
    assign memory[1297] = 12'h998;
    assign memory[1298] = 12'h998;
    assign memory[1299] = 12'h999;
    assign memory[1300] = 12'h998;
    assign memory[1301] = 12'h999;
    assign memory[1302] = 12'h999;
    assign memory[1303] = 12'h998;
    assign memory[1304] = 12'h999;
    assign memory[1305] = 12'h999;
    assign memory[1306] = 12'h998;
    assign memory[1307] = 12'h998;
    assign memory[1308] = 12'h898;
    assign memory[1309] = 12'h998;
    assign memory[1310] = 12'h998;
    assign memory[1311] = 12'h998;
    assign memory[1312] = 12'h998;
    assign memory[1313] = 12'h888;
    assign memory[1314] = 12'h999;
    assign memory[1315] = 12'h998;
    assign memory[1316] = 12'h888;
    assign memory[1317] = 12'h888;
    assign memory[1318] = 12'h898;
    assign memory[1319] = 12'h998;
    assign memory[1320] = 12'h898;
    assign memory[1321] = 12'h999;
    assign memory[1322] = 12'h998;
    assign memory[1323] = 12'h999;
    assign memory[1324] = 12'h888;
    assign memory[1325] = 12'h998;
    assign memory[1326] = 12'h888;
    assign memory[1327] = 12'h888;
    assign memory[1328] = 12'h998;
    assign memory[1329] = 12'h999;
    assign memory[1330] = 12'h999;
    assign memory[1331] = 12'h998;
    assign memory[1332] = 12'h998;
    assign memory[1333] = 12'h888;
    assign memory[1334] = 12'h998;
    assign memory[1335] = 12'h998;
    assign memory[1336] = 12'h888;
    assign memory[1337] = 12'h887;
    assign memory[1338] = 12'h998;
    assign memory[1339] = 12'h888;
    assign memory[1340] = 12'h998;
    assign memory[1341] = 12'h888;
    assign memory[1342] = 12'h998;
    assign memory[1343] = 12'h998;
    assign memory[1344] = 12'h999;
    assign memory[1345] = 12'h998;
    assign memory[1346] = 12'h888;
    assign memory[1347] = 12'h888;
    assign memory[1348] = 12'h888;
    assign memory[1349] = 12'h998;
    assign memory[1350] = 12'h998;
    assign memory[1351] = 12'h888;
    assign memory[1352] = 12'h998;
    assign memory[1353] = 12'h898;
    assign memory[1354] = 12'h888;
    assign memory[1355] = 12'h888;
    assign memory[1356] = 12'h998;
    assign memory[1357] = 12'h888;
    assign memory[1358] = 12'h998;
    assign memory[1359] = 12'h888;
    assign memory[1360] = 12'h999;
    assign memory[1361] = 12'h888;
    assign memory[1362] = 12'h998;
    assign memory[1363] = 12'h888;
    assign memory[1364] = 12'h998;
    assign memory[1365] = 12'h888;
    assign memory[1366] = 12'h888;
    assign memory[1367] = 12'h888;
    assign memory[1368] = 12'h998;
    assign memory[1369] = 12'h998;
    assign memory[1370] = 12'h998;
    assign memory[1371] = 12'h998;
    assign memory[1372] = 12'h998;
    assign memory[1373] = 12'h888;
    assign memory[1374] = 12'h998;
    assign memory[1375] = 12'h999;
    assign memory[1376] = 12'h888;
    assign memory[1377] = 12'h888;
    assign memory[1378] = 12'h998;
    assign memory[1379] = 12'h888;
    assign memory[1380] = 12'h999;
    assign memory[1381] = 12'h888;
    assign memory[1382] = 12'h998;
    assign memory[1383] = 12'h888;
    assign memory[1384] = 12'h888;
    assign memory[1385] = 12'h998;
    assign memory[1386] = 12'h999;
    assign memory[1387] = 12'h998;
    assign memory[1388] = 12'h999;
    assign memory[1389] = 12'h998;
    assign memory[1390] = 12'h999;
    assign memory[1391] = 12'h888;
    assign memory[1392] = 12'h898;
    assign memory[1393] = 12'h999;
    assign memory[1394] = 12'h998;
    assign memory[1395] = 12'h888;
    assign memory[1396] = 12'h998;
    assign memory[1397] = 12'h898;
    assign memory[1398] = 12'h999;
    assign memory[1399] = 12'h888;
    assign memory[1400] = 12'h998;
    assign memory[1401] = 12'h888;
    assign memory[1402] = 12'h898;
    assign memory[1403] = 12'h998;
    assign memory[1404] = 12'h888;
    assign memory[1405] = 12'h888;
    assign memory[1406] = 12'h887;
    assign memory[1407] = 12'h999;
    assign memory[1408] = 12'h998;
    assign memory[1409] = 12'h999;
    assign memory[1410] = 12'h888;
    assign memory[1411] = 12'h888;
    assign memory[1412] = 12'h998;
    assign memory[1413] = 12'h998;
    assign memory[1414] = 12'h888;
    assign memory[1415] = 12'h888;
    assign memory[1416] = 12'h998;
    assign memory[1417] = 12'h998;
    assign memory[1418] = 12'h898;
    assign memory[1419] = 12'h888;
    assign memory[1420] = 12'h888;
    assign memory[1421] = 12'h888;
    assign memory[1422] = 12'h887;
    assign memory[1423] = 12'h999;
    assign memory[1424] = 12'h888;
    assign memory[1425] = 12'h999;
    assign memory[1426] = 12'h888;
    assign memory[1427] = 12'h888;
    assign memory[1428] = 12'h999;
    assign memory[1429] = 12'h998;
    assign memory[1430] = 12'h998;
    assign memory[1431] = 12'h999;
    assign memory[1432] = 12'h999;
    assign memory[1433] = 12'h998;
    assign memory[1434] = 12'h999;
    assign memory[1435] = 12'h998;
    assign memory[1436] = 12'h998;
    assign memory[1437] = 12'h998;
    assign memory[1438] = 12'h998;
    assign memory[1439] = 12'h998;
    assign memory[1440] = 12'h998;
    assign memory[1441] = 12'h888;
    assign memory[1442] = 12'h998;
    assign memory[1443] = 12'h998;
    assign memory[1444] = 12'h998;
    assign memory[1445] = 12'h998;
    assign memory[1446] = 12'h998;
    assign memory[1447] = 12'h998;
    assign memory[1448] = 12'h998;
    assign memory[1449] = 12'h998;
    assign memory[1450] = 12'h888;
    assign memory[1451] = 12'h998;
    assign memory[1452] = 12'h999;
    assign memory[1453] = 12'h888;
    assign memory[1454] = 12'h998;
    assign memory[1455] = 12'h888;
    assign memory[1456] = 12'h998;
    assign memory[1457] = 12'h998;
    assign memory[1458] = 12'h998;
    assign memory[1459] = 12'h998;
    assign memory[1460] = 12'h888;
    assign memory[1461] = 12'h888;
    assign memory[1462] = 12'h998;
    assign memory[1463] = 12'h998;
    assign memory[1464] = 12'h998;
    assign memory[1465] = 12'h998;
    assign memory[1466] = 12'h998;
    assign memory[1467] = 12'h998;
    assign memory[1468] = 12'h888;
    assign memory[1469] = 12'h888;
    assign memory[1470] = 12'h999;
    assign memory[1471] = 12'h998;
    assign memory[1472] = 12'h998;
    assign memory[1473] = 12'h998;
    assign memory[1474] = 12'h898;
    assign memory[1475] = 12'h999;
    assign memory[1476] = 12'h888;
    assign memory[1477] = 12'h887;
    assign memory[1478] = 12'h998;
    assign memory[1479] = 12'h998;
    assign memory[1480] = 12'h998;
    assign memory[1481] = 12'h998;
    assign memory[1482] = 12'h998;
    assign memory[1483] = 12'h998;
    assign memory[1484] = 12'h998;
    assign memory[1485] = 12'h999;
    assign memory[1486] = 12'h888;
    assign memory[1487] = 12'h998;
    assign memory[1488] = 12'h998;
    assign memory[1489] = 12'h998;
    assign memory[1490] = 12'h998;
    assign memory[1491] = 12'h898;
    assign memory[1492] = 12'h888;
    assign memory[1493] = 12'h999;
    assign memory[1494] = 12'h888;
    assign memory[1495] = 12'h888;
    assign memory[1496] = 12'h999;
    assign memory[1497] = 12'h888;
    assign memory[1498] = 12'h898;
    assign memory[1499] = 12'h998;
    assign memory[1500] = 12'h999;
    assign memory[1501] = 12'h887;
    assign memory[1502] = 12'h998;
    assign memory[1503] = 12'h998;
    assign memory[1504] = 12'h887;
    assign memory[1505] = 12'h998;
    assign memory[1506] = 12'h888;
    assign memory[1507] = 12'h998;
    assign memory[1508] = 12'h888;
    assign memory[1509] = 12'h998;
    assign memory[1510] = 12'h998;
    assign memory[1511] = 12'h998;
    assign memory[1512] = 12'h888;
    assign memory[1513] = 12'h998;
    assign memory[1514] = 12'h998;
    assign memory[1515] = 12'h998;
    assign memory[1516] = 12'h998;
    assign memory[1517] = 12'h888;
    assign memory[1518] = 12'h898;
    assign memory[1519] = 12'h998;
    assign memory[1520] = 12'h888;
    assign memory[1521] = 12'h998;
    assign memory[1522] = 12'h998;
    assign memory[1523] = 12'h998;
    assign memory[1524] = 12'h888;
    assign memory[1525] = 12'h998;
    assign memory[1526] = 12'h888;
    assign memory[1527] = 12'h998;
    assign memory[1528] = 12'h888;
    assign memory[1529] = 12'h887;
    assign memory[1530] = 12'h888;
    assign memory[1531] = 12'h888;
    assign memory[1532] = 12'h888;
    assign memory[1533] = 12'h998;
    assign memory[1534] = 12'h998;
    assign memory[1535] = 12'h998;
    assign memory[1536] = 12'h998;
    assign memory[1537] = 12'h998;
    assign memory[1538] = 12'h998;
    assign memory[1539] = 12'h998;
    assign memory[1540] = 12'h998;
    assign memory[1541] = 12'h998;
    assign memory[1542] = 12'h998;
    assign memory[1543] = 12'h998;
    assign memory[1544] = 12'h888;
    assign memory[1545] = 12'h888;
    assign memory[1546] = 12'h998;
    assign memory[1547] = 12'h888;
    assign memory[1548] = 12'h888;
    assign memory[1549] = 12'h998;
    assign memory[1550] = 12'h998;
    assign memory[1551] = 12'h998;
    assign memory[1552] = 12'h998;
    assign memory[1553] = 12'h998;
    assign memory[1554] = 12'h888;
    assign memory[1555] = 12'h998;
    assign memory[1556] = 12'h998;
    assign memory[1557] = 12'h998;
    assign memory[1558] = 12'h998;
    assign memory[1559] = 12'h888;
    assign memory[1560] = 12'h998;
    assign memory[1561] = 12'h998;
    assign memory[1562] = 12'h998;
    assign memory[1563] = 12'h998;
    assign memory[1564] = 12'h998;
    assign memory[1565] = 12'h888;
    assign memory[1566] = 12'h998;
    assign memory[1567] = 12'h887;
    assign memory[1568] = 12'h888;
    assign memory[1569] = 12'h888;
    assign memory[1570] = 12'h998;
    assign memory[1571] = 12'h999;
    assign memory[1572] = 12'h999;
    assign memory[1573] = 12'h888;
    assign memory[1574] = 12'h998;
    assign memory[1575] = 12'h998;
    assign memory[1576] = 12'h898;
    assign memory[1577] = 12'h998;
    assign memory[1578] = 12'h999;
    assign memory[1579] = 12'h998;
    assign memory[1580] = 12'h888;
    assign memory[1581] = 12'h888;
    assign memory[1582] = 12'h998;
    assign memory[1583] = 12'h998;
    assign memory[1584] = 12'h998;
    assign memory[1585] = 12'h898;
    assign memory[1586] = 12'h998;
    assign memory[1587] = 12'h998;
    assign memory[1588] = 12'h998;
    assign memory[1589] = 12'h998;
    assign memory[1590] = 12'h998;
    assign memory[1591] = 12'h998;
    assign memory[1592] = 12'h998;
    assign memory[1593] = 12'h999;
    assign memory[1594] = 12'h999;
    assign memory[1595] = 12'h998;
    assign memory[1596] = 12'h888;
    assign memory[1597] = 12'h998;
    assign memory[1598] = 12'h998;
    assign memory[1599] = 12'h998;
    assign memory[1600] = 12'h999;
    assign memory[1601] = 12'h998;
    assign memory[1602] = 12'h999;
    assign memory[1603] = 12'h888;
    assign memory[1604] = 12'h999;
    assign memory[1605] = 12'h888;
    assign memory[1606] = 12'h998;
    assign memory[1607] = 12'h998;
    assign memory[1608] = 12'h998;
    assign memory[1609] = 12'h998;
    assign memory[1610] = 12'h998;
    assign memory[1611] = 12'h888;
    assign memory[1612] = 12'h998;
    assign memory[1613] = 12'h999;
    assign memory[1614] = 12'h999;
    assign memory[1615] = 12'h999;
    assign memory[1616] = 12'h998;
    assign memory[1617] = 12'h999;
    assign memory[1618] = 12'h998;
    assign memory[1619] = 12'h999;
    assign memory[1620] = 12'h888;
    assign memory[1621] = 12'h998;
    assign memory[1622] = 12'h998;
    assign memory[1623] = 12'h998;
    assign memory[1624] = 12'h888;
    assign memory[1625] = 12'h999;
    assign memory[1626] = 12'h998;
    assign memory[1627] = 12'h888;
    assign memory[1628] = 12'h888;
    assign memory[1629] = 12'h998;
    assign memory[1630] = 12'h998;
    assign memory[1631] = 12'h999;
    assign memory[1632] = 12'h999;
    assign memory[1633] = 12'h998;
    assign memory[1634] = 12'h888;
    assign memory[1635] = 12'h998;
    assign memory[1636] = 12'h999;
    assign memory[1637] = 12'h999;
    assign memory[1638] = 12'h998;
    assign memory[1639] = 12'h998;
    assign memory[1640] = 12'h998;
    assign memory[1641] = 12'h888;
    assign memory[1642] = 12'h888;
    assign memory[1643] = 12'h998;
    assign memory[1644] = 12'h888;
    assign memory[1645] = 12'h898;
    assign memory[1646] = 12'h898;
    assign memory[1647] = 12'h888;
    assign memory[1648] = 12'h998;
    assign memory[1649] = 12'h998;
    assign memory[1650] = 12'h998;
    assign memory[1651] = 12'h998;
    assign memory[1652] = 12'h998;
    assign memory[1653] = 12'h998;
    assign memory[1654] = 12'h998;
    assign memory[1655] = 12'h998;
    assign memory[1656] = 12'h888;
    assign memory[1657] = 12'h888;
    assign memory[1658] = 12'h898;
    assign memory[1659] = 12'h998;
    assign memory[1660] = 12'h998;
    assign memory[1661] = 12'h998;
    assign memory[1662] = 12'h998;
    assign memory[1663] = 12'h888;
    assign memory[1664] = 12'h887;
    assign memory[1665] = 12'h999;
    assign memory[1666] = 12'h998;
    assign memory[1667] = 12'h888;
    assign memory[1668] = 12'h998;
    assign memory[1669] = 12'h998;
    assign memory[1670] = 12'h998;
    assign memory[1671] = 12'h898;
    assign memory[1672] = 12'h998;
    assign memory[1673] = 12'h998;
    assign memory[1674] = 12'h998;
    assign memory[1675] = 12'h998;
    assign memory[1676] = 12'h998;
    assign memory[1677] = 12'h888;
    assign memory[1678] = 12'h998;
    assign memory[1679] = 12'h998;
    assign memory[1680] = 12'h998;
    assign memory[1681] = 12'h999;
    assign memory[1682] = 12'h998;
    assign memory[1683] = 12'h998;
    assign memory[1684] = 12'h898;
    assign memory[1685] = 12'h999;
    assign memory[1686] = 12'h998;
    assign memory[1687] = 12'h998;
    assign memory[1688] = 12'h888;
    assign memory[1689] = 12'h998;
    assign memory[1690] = 12'h998;
    assign memory[1691] = 12'h999;
    assign memory[1692] = 12'h998;
    assign memory[1693] = 12'h998;
    assign memory[1694] = 12'h888;
    assign memory[1695] = 12'h888;
    assign memory[1696] = 12'h999;
    assign memory[1697] = 12'h999;
    assign memory[1698] = 12'h998;
    assign memory[1699] = 12'h999;
    assign memory[1700] = 12'h998;
    assign memory[1701] = 12'h888;
    assign memory[1702] = 12'h898;
    assign memory[1703] = 12'h999;
    assign memory[1704] = 12'h888;
    assign memory[1705] = 12'h888;
    assign memory[1706] = 12'h999;
    assign memory[1707] = 12'h998;
    assign memory[1708] = 12'h998;
    assign memory[1709] = 12'h999;
    assign memory[1710] = 12'h998;
    assign memory[1711] = 12'h998;
    assign memory[1712] = 12'h998;
    assign memory[1713] = 12'h898;
    assign memory[1714] = 12'h998;
    assign memory[1715] = 12'h998;
    assign memory[1716] = 12'h998;
    assign memory[1717] = 12'h998;
    assign memory[1718] = 12'h888;
    assign memory[1719] = 12'h999;
    assign memory[1720] = 12'h998;
    assign memory[1721] = 12'h888;
    assign memory[1722] = 12'h998;
    assign memory[1723] = 12'h888;
    assign memory[1724] = 12'h999;
    assign memory[1725] = 12'h998;
    assign memory[1726] = 12'h888;
    assign memory[1727] = 12'h888;
    assign memory[1728] = 12'h998;
    assign memory[1729] = 12'h998;
    assign memory[1730] = 12'h999;
    assign memory[1731] = 12'h998;
    assign memory[1732] = 12'h999;
    assign memory[1733] = 12'h888;
    assign memory[1734] = 12'h999;
    assign memory[1735] = 12'h888;
    assign memory[1736] = 12'h998;
    assign memory[1737] = 12'h998;
    assign memory[1738] = 12'h998;
    assign memory[1739] = 12'h998;
    assign memory[1740] = 12'h998;
    assign memory[1741] = 12'h888;
    assign memory[1742] = 12'h998;
    assign memory[1743] = 12'h999;
    assign memory[1744] = 12'h999;
    assign memory[1745] = 12'h999;
    assign memory[1746] = 12'h998;
    assign memory[1747] = 12'h999;
    assign memory[1748] = 12'h998;
    assign memory[1749] = 12'h999;
    assign memory[1750] = 12'h888;
    assign memory[1751] = 12'h998;
    assign memory[1752] = 12'h998;
    assign memory[1753] = 12'h998;
    assign memory[1754] = 12'h888;
    assign memory[1755] = 12'h999;
    assign memory[1756] = 12'h998;
    assign memory[1757] = 12'h888;
    assign memory[1758] = 12'h888;
    assign memory[1759] = 12'h998;
    assign memory[1760] = 12'h998;
    assign memory[1761] = 12'h998;
    assign memory[1762] = 12'h998;
    assign memory[1763] = 12'h998;
    assign memory[1764] = 12'h998;
    assign memory[1765] = 12'h898;
    assign memory[1766] = 12'h998;
    assign memory[1767] = 12'h998;
    assign memory[1768] = 12'h998;
    assign memory[1769] = 12'h998;
    assign memory[1770] = 12'h999;
    assign memory[1771] = 12'h888;
    assign memory[1772] = 12'h898;
    assign memory[1773] = 12'h888;
    assign memory[1774] = 12'h998;
    assign memory[1775] = 12'h999;
    assign memory[1776] = 12'h998;
    assign memory[1777] = 12'h898;
    assign memory[1778] = 12'h999;
    assign memory[1779] = 12'h998;
    assign memory[1780] = 12'h998;
    assign memory[1781] = 12'h998;
    assign memory[1782] = 12'h998;
    assign memory[1783] = 12'h999;
    assign memory[1784] = 12'h998;
    assign memory[1785] = 12'h888;
    assign memory[1786] = 12'h888;
    assign memory[1787] = 12'h888;
    assign memory[1788] = 12'h898;
    assign memory[1789] = 12'h999;
    assign memory[1790] = 12'h998;
    assign memory[1791] = 12'h888;
    assign memory[1792] = 12'h888;
    assign memory[1793] = 12'h998;
    assign memory[1794] = 12'h888;
    assign memory[1795] = 12'h888;
    assign memory[1796] = 12'h998;
    assign memory[1797] = 12'h888;
    assign memory[1798] = 12'h998;
    assign memory[1799] = 12'h888;
    assign memory[1800] = 12'h998;
    assign memory[1801] = 12'h999;
    assign memory[1802] = 12'h888;
    assign memory[1803] = 12'h998;
    assign memory[1804] = 12'h898;
    assign memory[1805] = 12'h998;
    assign memory[1806] = 12'h888;
    assign memory[1807] = 12'h887;
    assign memory[1808] = 12'h998;
    assign memory[1809] = 12'h999;
    assign memory[1810] = 12'h999;
    assign memory[1811] = 12'h888;
    assign memory[1812] = 12'h998;
    assign memory[1813] = 12'h888;
    assign memory[1814] = 12'h998;
    assign memory[1815] = 12'h888;
    assign memory[1816] = 12'h998;
    assign memory[1817] = 12'h998;
    assign memory[1818] = 12'h999;
    assign memory[1819] = 12'h888;
    assign memory[1820] = 12'h888;
    assign memory[1821] = 12'h998;
    assign memory[1822] = 12'h888;
    assign memory[1823] = 12'h999;
    assign memory[1824] = 12'h888;
    assign memory[1825] = 12'h888;
    assign memory[1826] = 12'h998;
    assign memory[1827] = 12'h998;
    assign memory[1828] = 12'h898;
    assign memory[1829] = 12'h998;
    assign memory[1830] = 12'h998;
    assign memory[1831] = 12'h998;
    assign memory[1832] = 12'h888;
    assign memory[1833] = 12'h888;
    assign memory[1834] = 12'h998;
    assign memory[1835] = 12'h888;
    assign memory[1836] = 12'h888;
    assign memory[1837] = 12'h998;
    assign memory[1838] = 12'h888;
    assign memory[1839] = 12'h998;
    assign memory[1840] = 12'h888;
    assign memory[1841] = 12'h998;
    assign memory[1842] = 12'h998;
    assign memory[1843] = 12'h888;
    assign memory[1844] = 12'h998;
    assign memory[1845] = 12'h999;
    assign memory[1846] = 12'h888;
    assign memory[1847] = 12'h998;
    assign memory[1848] = 12'h998;
    assign memory[1849] = 12'h998;
    assign memory[1850] = 12'h998;
    assign memory[1851] = 12'h998;
    assign memory[1852] = 12'h888;
    assign memory[1853] = 12'h888;
    assign memory[1854] = 12'h998;
    assign memory[1855] = 12'h999;
    assign memory[1856] = 12'h998;
    assign memory[1857] = 12'h998;
    assign memory[1858] = 12'h998;
    assign memory[1859] = 12'h998;
    assign memory[1860] = 12'h998;
    assign memory[1861] = 12'h998;
    assign memory[1862] = 12'h998;
    assign memory[1863] = 12'h998;
    assign memory[1864] = 12'h998;
    assign memory[1865] = 12'h898;
    assign memory[1866] = 12'h898;
    assign memory[1867] = 12'h998;
    assign memory[1868] = 12'h888;
    assign memory[1869] = 12'h998;
    assign memory[1870] = 12'h998;
    assign memory[1871] = 12'h998;
    assign memory[1872] = 12'h998;
    assign memory[1873] = 12'h998;
    assign memory[1874] = 12'h999;
    assign memory[1875] = 12'h998;
    assign memory[1876] = 12'h998;
    assign memory[1877] = 12'h998;
    assign memory[1878] = 12'h998;
    assign memory[1879] = 12'h999;
    assign memory[1880] = 12'h888;
    assign memory[1881] = 12'h998;
    assign memory[1882] = 12'h887;
    assign memory[1883] = 12'h888;
    assign memory[1884] = 12'h998;
    assign memory[1885] = 12'h998;
    assign memory[1886] = 12'h998;
    assign memory[1887] = 12'h898;
    assign memory[1888] = 12'h999;
    assign memory[1889] = 12'h999;
    assign memory[1890] = 12'h998;
    assign memory[1891] = 12'h888;
    assign memory[1892] = 12'h998;
    assign memory[1893] = 12'h998;
    assign memory[1894] = 12'h998;
    assign memory[1895] = 12'h888;
    assign memory[1896] = 12'h998;
    assign memory[1897] = 12'h998;
    assign memory[1898] = 12'h887;
    assign memory[1899] = 12'h888;
    assign memory[1900] = 12'h888;
    assign memory[1901] = 12'h999;
    assign memory[1902] = 12'h888;
    assign memory[1903] = 12'h999;
    assign memory[1904] = 12'h998;
    assign memory[1905] = 12'h999;
    assign memory[1906] = 12'h888;
    assign memory[1907] = 12'h998;
    assign memory[1908] = 12'h998;
    assign memory[1909] = 12'h998;
    assign memory[1910] = 12'h898;
    assign memory[1911] = 12'h998;
    assign memory[1912] = 12'h999;
    assign memory[1913] = 12'h998;
    assign memory[1914] = 12'h888;
    assign memory[1915] = 12'h998;
    assign memory[1916] = 12'h888;
    assign memory[1917] = 12'h998;
    assign memory[1918] = 12'h998;
    assign memory[1919] = 12'h998;
    assign memory[1920] = 12'h888;
    assign memory[1921] = 12'h999;
    assign memory[1922] = 12'h998;
    assign memory[1923] = 12'h888;
    assign memory[1924] = 12'h898;
    assign memory[1925] = 12'h998;
    assign memory[1926] = 12'h898;
    assign memory[1927] = 12'h998;
    assign memory[1928] = 12'h998;
    assign memory[1929] = 12'h998;
    assign memory[1930] = 12'h888;
    assign memory[1931] = 12'h999;
    assign memory[1932] = 12'h888;
    assign memory[1933] = 12'h998;
    assign memory[1934] = 12'h998;
    assign memory[1935] = 12'h999;
    assign memory[1936] = 12'h998;
    assign memory[1937] = 12'h888;
    assign memory[1938] = 12'h998;
    assign memory[1939] = 12'h888;
    assign memory[1940] = 12'h998;
    assign memory[1941] = 12'h888;
    assign memory[1942] = 12'h888;
    assign memory[1943] = 12'h999;
    assign memory[1944] = 12'h998;
    assign memory[1945] = 12'h887;
    assign memory[1946] = 12'h999;
    assign memory[1947] = 12'h998;
    assign memory[1948] = 12'h998;
    assign memory[1949] = 12'h998;
    assign memory[1950] = 12'h888;
    assign memory[1951] = 12'h998;
    assign memory[1952] = 12'h998;
    assign memory[1953] = 12'h998;
    assign memory[1954] = 12'h888;
    assign memory[1955] = 12'h888;
    assign memory[1956] = 12'h998;
    assign memory[1957] = 12'h888;
    assign memory[1958] = 12'h888;
    assign memory[1959] = 12'h998;
    assign memory[1960] = 12'h998;
    assign memory[1961] = 12'h998;
    assign memory[1962] = 12'h998;
    assign memory[1963] = 12'h998;
    assign memory[1964] = 12'h888;
    assign memory[1965] = 12'h998;
    assign memory[1966] = 12'h998;
    assign memory[1967] = 12'h998;
    assign memory[1968] = 12'h998;
    assign memory[1969] = 12'h888;
    assign memory[1970] = 12'h998;
    assign memory[1971] = 12'h998;
    assign memory[1972] = 12'h998;
    assign memory[1973] = 12'h998;
    assign memory[1974] = 12'h998;
    assign memory[1975] = 12'h888;
    assign memory[1976] = 12'h998;
    assign memory[1977] = 12'h887;
    assign memory[1978] = 12'h998;
    assign memory[1979] = 12'h998;
    assign memory[1980] = 12'h998;
    assign memory[1981] = 12'h998;
    assign memory[1982] = 12'h998;
    assign memory[1983] = 12'h998;
    assign memory[1984] = 12'h998;
    assign memory[1985] = 12'h998;
    assign memory[1986] = 12'h999;
    assign memory[1987] = 12'h999;
    assign memory[1988] = 12'h998;
    assign memory[1989] = 12'h999;
    assign memory[1990] = 12'h998;
    assign memory[1991] = 12'h998;
    assign memory[1992] = 12'h998;
    assign memory[1993] = 12'h888;
    assign memory[1994] = 12'h888;
    assign memory[1995] = 12'h998;
    assign memory[1996] = 12'h998;
    assign memory[1997] = 12'h898;
    assign memory[1998] = 12'h898;
    assign memory[1999] = 12'h998;
    assign memory[2000] = 12'h998;
    assign memory[2001] = 12'h998;
    assign memory[2002] = 12'h998;
    assign memory[2003] = 12'h999;
    assign memory[2004] = 12'h888;
    assign memory[2005] = 12'h888;
    assign memory[2006] = 12'h998;
    assign memory[2007] = 12'h998;
    assign memory[2008] = 12'h998;
    assign memory[2009] = 12'h998;
    assign memory[2010] = 12'h998;
    assign memory[2011] = 12'h998;
    assign memory[2012] = 12'h998;
    assign memory[2013] = 12'h998;
    assign memory[2014] = 12'h998;
    assign memory[2015] = 12'h888;
    assign memory[2016] = 12'h888;
    assign memory[2017] = 12'h888;
    assign memory[2018] = 12'h998;
    assign memory[2019] = 12'h998;
    assign memory[2020] = 12'h999;
    assign memory[2021] = 12'h998;
    assign memory[2022] = 12'h888;
    assign memory[2023] = 12'h998;
    assign memory[2024] = 12'h888;
    assign memory[2025] = 12'h999;
    assign memory[2026] = 12'h888;
    assign memory[2027] = 12'h888;
    assign memory[2028] = 12'h999;
    assign memory[2029] = 12'h999;
    assign memory[2030] = 12'h998;
    assign memory[2031] = 12'h888;
    assign memory[2032] = 12'h998;
    assign memory[2033] = 12'h998;
    assign memory[2034] = 12'h999;
    assign memory[2035] = 12'h998;
    assign memory[2036] = 12'h888;
    assign memory[2037] = 12'h998;
    assign memory[2038] = 12'h898;
    assign memory[2039] = 12'h887;
    assign memory[2040] = 12'h998;
    assign memory[2041] = 12'h888;
    assign memory[2042] = 12'h998;
    assign memory[2043] = 12'h888;
    assign memory[2044] = 12'h998;
    assign memory[2045] = 12'h998;
    assign memory[2046] = 12'h998;
    assign memory[2047] = 12'h998;
    assign memory[2048] = 12'h000;
    assign memory[2049] = 12'h000;
    assign memory[2050] = 12'h000;
    assign memory[2051] = 12'h000;
    assign memory[2052] = 12'h000;
    assign memory[2053] = 12'h000;
    assign memory[2054] = 12'h000;
    assign memory[2055] = 12'h000;
    assign memory[2056] = 12'h000;
    assign memory[2057] = 12'h000;
    assign memory[2058] = 12'h000;
    assign memory[2059] = 12'h000;
    assign memory[2060] = 12'h000;
    assign memory[2061] = 12'h000;
    assign memory[2062] = 12'h000;
    assign memory[2063] = 12'h000;
    assign memory[2064] = 12'h000;
    assign memory[2065] = 12'h000;
    assign memory[2066] = 12'h000;
    assign memory[2067] = 12'h000;
    assign memory[2068] = 12'h000;
    assign memory[2069] = 12'h000;
    assign memory[2070] = 12'h000;
    assign memory[2071] = 12'h000;
    assign memory[2072] = 12'h000;
    assign memory[2073] = 12'h000;
    assign memory[2074] = 12'h000;
    assign memory[2075] = 12'h000;
    assign memory[2076] = 12'h000;
    assign memory[2077] = 12'h000;
    assign memory[2078] = 12'h000;
    assign memory[2079] = 12'h000;
    assign memory[2080] = 12'h000;
    assign memory[2081] = 12'h000;
    assign memory[2082] = 12'h000;
    assign memory[2083] = 12'h000;
    assign memory[2084] = 12'h000;
    assign memory[2085] = 12'h000;
    assign memory[2086] = 12'h000;
    assign memory[2087] = 12'h000;
    assign memory[2088] = 12'h000;
    assign memory[2089] = 12'h000;
    assign memory[2090] = 12'h000;
    assign memory[2091] = 12'h000;
    assign memory[2092] = 12'h000;
    assign memory[2093] = 12'h000;
    assign memory[2094] = 12'h000;
    assign memory[2095] = 12'h000;
    assign memory[2096] = 12'h000;
    assign memory[2097] = 12'h000;
    assign memory[2098] = 12'h000;
    assign memory[2099] = 12'h000;
    assign memory[2100] = 12'h000;
    assign memory[2101] = 12'h000;
    assign memory[2102] = 12'h000;
    assign memory[2103] = 12'h000;
    assign memory[2104] = 12'h000;
    assign memory[2105] = 12'h000;
    assign memory[2106] = 12'h000;
    assign memory[2107] = 12'h000;
    assign memory[2108] = 12'h000;
    assign memory[2109] = 12'h000;
    assign memory[2110] = 12'h000;
    assign memory[2111] = 12'h000;
    assign memory[2112] = 12'h000;
    assign memory[2113] = 12'h000;
    assign memory[2114] = 12'h000;
    assign memory[2115] = 12'h000;
    assign memory[2116] = 12'h000;
    assign memory[2117] = 12'h000;
    assign memory[2118] = 12'h000;
    assign memory[2119] = 12'h000;
    assign memory[2120] = 12'h000;
    assign memory[2121] = 12'h000;
    assign memory[2122] = 12'h000;
    assign memory[2123] = 12'h000;
    assign memory[2124] = 12'h000;
    assign memory[2125] = 12'h000;
    assign memory[2126] = 12'h000;
    assign memory[2127] = 12'h000;
    assign memory[2128] = 12'h000;
    assign memory[2129] = 12'h000;
    assign memory[2130] = 12'h000;
    assign memory[2131] = 12'h000;
    assign memory[2132] = 12'h000;
    assign memory[2133] = 12'h000;
    assign memory[2134] = 12'h000;
    assign memory[2135] = 12'h000;
    assign memory[2136] = 12'h000;
    assign memory[2137] = 12'h000;
    assign memory[2138] = 12'h000;
    assign memory[2139] = 12'h000;
    assign memory[2140] = 12'h000;
    assign memory[2141] = 12'h000;
    assign memory[2142] = 12'h000;
    assign memory[2143] = 12'h000;
    assign memory[2144] = 12'h000;
    assign memory[2145] = 12'h000;
    assign memory[2146] = 12'h000;
    assign memory[2147] = 12'h000;
    assign memory[2148] = 12'h000;
    assign memory[2149] = 12'h000;
    assign memory[2150] = 12'h000;
    assign memory[2151] = 12'h000;
    assign memory[2152] = 12'h000;
    assign memory[2153] = 12'h000;
    assign memory[2154] = 12'h000;
    assign memory[2155] = 12'h000;
    assign memory[2156] = 12'h000;
    assign memory[2157] = 12'h000;
    assign memory[2158] = 12'h000;
    assign memory[2159] = 12'h000;
    assign memory[2160] = 12'h000;
    assign memory[2161] = 12'h000;
    assign memory[2162] = 12'h000;
    assign memory[2163] = 12'h000;
    assign memory[2164] = 12'h000;
    assign memory[2165] = 12'h000;
    assign memory[2166] = 12'h000;
    assign memory[2167] = 12'h000;
    assign memory[2168] = 12'h000;
    assign memory[2169] = 12'h000;
    assign memory[2170] = 12'h000;
    assign memory[2171] = 12'h000;
    assign memory[2172] = 12'h000;
    assign memory[2173] = 12'h000;
    assign memory[2174] = 12'h000;
    assign memory[2175] = 12'h000;
    assign memory[2176] = 12'h000;
    assign memory[2177] = 12'h000;
    assign memory[2178] = 12'h000;
    assign memory[2179] = 12'h000;
    assign memory[2180] = 12'h000;
    assign memory[2181] = 12'h000;
    assign memory[2182] = 12'h000;
    assign memory[2183] = 12'h000;
    assign memory[2184] = 12'h000;
    assign memory[2185] = 12'h000;
    assign memory[2186] = 12'h000;
    assign memory[2187] = 12'h000;
    assign memory[2188] = 12'h000;
    assign memory[2189] = 12'h000;
    assign memory[2190] = 12'h000;
    assign memory[2191] = 12'h000;
    assign memory[2192] = 12'h000;
    assign memory[2193] = 12'h000;
    assign memory[2194] = 12'h000;
    assign memory[2195] = 12'h000;
    assign memory[2196] = 12'h000;
    assign memory[2197] = 12'h000;
    assign memory[2198] = 12'h000;
    assign memory[2199] = 12'h000;
    assign memory[2200] = 12'h000;
    assign memory[2201] = 12'h000;
    assign memory[2202] = 12'h000;
    assign memory[2203] = 12'h000;
    assign memory[2204] = 12'h000;
    assign memory[2205] = 12'h000;
    assign memory[2206] = 12'h000;
    assign memory[2207] = 12'h000;
    assign memory[2208] = 12'h000;
    assign memory[2209] = 12'h000;
    assign memory[2210] = 12'h000;
    assign memory[2211] = 12'h000;
    assign memory[2212] = 12'h000;
    assign memory[2213] = 12'h000;
    assign memory[2214] = 12'h000;
    assign memory[2215] = 12'h000;
    assign memory[2216] = 12'h000;
    assign memory[2217] = 12'h000;
    assign memory[2218] = 12'h000;
    assign memory[2219] = 12'h000;
    assign memory[2220] = 12'h000;
    assign memory[2221] = 12'h000;
    assign memory[2222] = 12'h000;
    assign memory[2223] = 12'h000;
    assign memory[2224] = 12'h000;
    assign memory[2225] = 12'h000;
    assign memory[2226] = 12'h000;
    assign memory[2227] = 12'h000;
    assign memory[2228] = 12'h000;
    assign memory[2229] = 12'h000;
    assign memory[2230] = 12'h000;
    assign memory[2231] = 12'h000;
    assign memory[2232] = 12'h000;
    assign memory[2233] = 12'h000;
    assign memory[2234] = 12'h000;
    assign memory[2235] = 12'h000;
    assign memory[2236] = 12'h000;
    assign memory[2237] = 12'h000;
    assign memory[2238] = 12'h000;
    assign memory[2239] = 12'h000;
    assign memory[2240] = 12'h000;
    assign memory[2241] = 12'h000;
    assign memory[2242] = 12'h000;
    assign memory[2243] = 12'h000;
    assign memory[2244] = 12'h000;
    assign memory[2245] = 12'h000;
    assign memory[2246] = 12'h000;
    assign memory[2247] = 12'h000;
    assign memory[2248] = 12'h000;
    assign memory[2249] = 12'h000;
    assign memory[2250] = 12'h000;
    assign memory[2251] = 12'h000;
    assign memory[2252] = 12'h000;
    assign memory[2253] = 12'h000;
    assign memory[2254] = 12'h000;
    assign memory[2255] = 12'h000;
    assign memory[2256] = 12'h000;
    assign memory[2257] = 12'h000;
    assign memory[2258] = 12'h000;
    assign memory[2259] = 12'h000;
    assign memory[2260] = 12'h000;
    assign memory[2261] = 12'h000;
    assign memory[2262] = 12'h000;
    assign memory[2263] = 12'h000;
    assign memory[2264] = 12'h000;
    assign memory[2265] = 12'h000;
    assign memory[2266] = 12'h000;
    assign memory[2267] = 12'h000;
    assign memory[2268] = 12'h000;
    assign memory[2269] = 12'h000;
    assign memory[2270] = 12'h000;
    assign memory[2271] = 12'h000;
    assign memory[2272] = 12'h000;
    assign memory[2273] = 12'h000;
    assign memory[2274] = 12'h000;
    assign memory[2275] = 12'h000;
    assign memory[2276] = 12'h000;
    assign memory[2277] = 12'h000;
    assign memory[2278] = 12'h000;
    assign memory[2279] = 12'h000;
    assign memory[2280] = 12'h000;
    assign memory[2281] = 12'h000;
    assign memory[2282] = 12'h000;
    assign memory[2283] = 12'h000;
    assign memory[2284] = 12'h000;
    assign memory[2285] = 12'h000;
    assign memory[2286] = 12'h000;
    assign memory[2287] = 12'h000;
    assign memory[2288] = 12'h000;
    assign memory[2289] = 12'h000;
    assign memory[2290] = 12'h000;
    assign memory[2291] = 12'h000;
    assign memory[2292] = 12'h000;
    assign memory[2293] = 12'h000;
    assign memory[2294] = 12'h000;
    assign memory[2295] = 12'h000;
    assign memory[2296] = 12'h000;
    assign memory[2297] = 12'h000;
    assign memory[2298] = 12'h000;
    assign memory[2299] = 12'h000;
    assign memory[2300] = 12'h000;
    assign memory[2301] = 12'h000;
    assign memory[2302] = 12'h000;
    assign memory[2303] = 12'h000;
    assign memory[2304] = 12'h000;
    assign memory[2305] = 12'h000;
    assign memory[2306] = 12'h000;
    assign memory[2307] = 12'h000;
    assign memory[2308] = 12'h000;
    assign memory[2309] = 12'h000;
    assign memory[2310] = 12'h000;
    assign memory[2311] = 12'h000;
    assign memory[2312] = 12'h000;
    assign memory[2313] = 12'h000;
    assign memory[2314] = 12'h000;
    assign memory[2315] = 12'h000;
    assign memory[2316] = 12'h000;
    assign memory[2317] = 12'h000;
    assign memory[2318] = 12'h000;
    assign memory[2319] = 12'h000;
    assign memory[2320] = 12'h000;
    assign memory[2321] = 12'h000;
    assign memory[2322] = 12'h000;
    assign memory[2323] = 12'h000;
    assign memory[2324] = 12'h000;
    assign memory[2325] = 12'h000;
    assign memory[2326] = 12'h000;
    assign memory[2327] = 12'h000;
    assign memory[2328] = 12'h000;
    assign memory[2329] = 12'h000;
    assign memory[2330] = 12'h000;
    assign memory[2331] = 12'h000;
    assign memory[2332] = 12'h000;
    assign memory[2333] = 12'h000;
    assign memory[2334] = 12'h000;
    assign memory[2335] = 12'h000;
    assign memory[2336] = 12'h000;
    assign memory[2337] = 12'h000;
    assign memory[2338] = 12'h000;
    assign memory[2339] = 12'h000;
    assign memory[2340] = 12'h000;
    assign memory[2341] = 12'h000;
    assign memory[2342] = 12'h000;
    assign memory[2343] = 12'h000;
    assign memory[2344] = 12'h000;
    assign memory[2345] = 12'h000;
    assign memory[2346] = 12'h000;
    assign memory[2347] = 12'h000;
    assign memory[2348] = 12'h000;
    assign memory[2349] = 12'h000;
    assign memory[2350] = 12'h000;
    assign memory[2351] = 12'h000;
    assign memory[2352] = 12'h000;
    assign memory[2353] = 12'h000;
    assign memory[2354] = 12'h000;
    assign memory[2355] = 12'h000;
    assign memory[2356] = 12'h000;
    assign memory[2357] = 12'h000;
    assign memory[2358] = 12'h000;
    assign memory[2359] = 12'h000;
    assign memory[2360] = 12'h000;
    assign memory[2361] = 12'h000;
    assign memory[2362] = 12'h000;
    assign memory[2363] = 12'h000;
    assign memory[2364] = 12'h000;
    assign memory[2365] = 12'h000;
    assign memory[2366] = 12'h000;
    assign memory[2367] = 12'h000;
    assign memory[2368] = 12'h000;
    assign memory[2369] = 12'h000;
    assign memory[2370] = 12'h000;
    assign memory[2371] = 12'h000;
    assign memory[2372] = 12'h000;
    assign memory[2373] = 12'h000;
    assign memory[2374] = 12'h000;
    assign memory[2375] = 12'h000;
    assign memory[2376] = 12'h000;
    assign memory[2377] = 12'h000;
    assign memory[2378] = 12'h000;
    assign memory[2379] = 12'h000;
    assign memory[2380] = 12'h000;
    assign memory[2381] = 12'h000;
    assign memory[2382] = 12'h000;
    assign memory[2383] = 12'h000;
    assign memory[2384] = 12'h000;
    assign memory[2385] = 12'h000;
    assign memory[2386] = 12'h000;
    assign memory[2387] = 12'h000;
    assign memory[2388] = 12'h000;
    assign memory[2389] = 12'h000;
    assign memory[2390] = 12'h000;
    assign memory[2391] = 12'h000;
    assign memory[2392] = 12'h000;
    assign memory[2393] = 12'h000;
    assign memory[2394] = 12'h000;
    assign memory[2395] = 12'h000;
    assign memory[2396] = 12'h000;
    assign memory[2397] = 12'h000;
    assign memory[2398] = 12'h000;
    assign memory[2399] = 12'h000;
    assign memory[2400] = 12'h000;
    assign memory[2401] = 12'h000;
    assign memory[2402] = 12'h000;
    assign memory[2403] = 12'h000;
    assign memory[2404] = 12'h000;
    assign memory[2405] = 12'h000;
    assign memory[2406] = 12'h000;
    assign memory[2407] = 12'h000;
    assign memory[2408] = 12'h000;
    assign memory[2409] = 12'h000;
    assign memory[2410] = 12'h000;
    assign memory[2411] = 12'h000;
    assign memory[2412] = 12'h000;
    assign memory[2413] = 12'h000;
    assign memory[2414] = 12'h000;
    assign memory[2415] = 12'h000;
    assign memory[2416] = 12'h000;
    assign memory[2417] = 12'h000;
    assign memory[2418] = 12'h000;
    assign memory[2419] = 12'h000;
    assign memory[2420] = 12'h000;
    assign memory[2421] = 12'h000;
    assign memory[2422] = 12'h000;
    assign memory[2423] = 12'h000;
    assign memory[2424] = 12'h000;
    assign memory[2425] = 12'h000;
    assign memory[2426] = 12'h000;
    assign memory[2427] = 12'h000;
    assign memory[2428] = 12'h000;
    assign memory[2429] = 12'h000;
    assign memory[2430] = 12'h000;
    assign memory[2431] = 12'h000;
    assign memory[2432] = 12'h000;
    assign memory[2433] = 12'h000;
    assign memory[2434] = 12'h000;
    assign memory[2435] = 12'h000;
    assign memory[2436] = 12'h000;
    assign memory[2437] = 12'h000;
    assign memory[2438] = 12'h000;
    assign memory[2439] = 12'h000;
    assign memory[2440] = 12'h000;
    assign memory[2441] = 12'h000;
    assign memory[2442] = 12'h000;
    assign memory[2443] = 12'h000;
    assign memory[2444] = 12'h000;
    assign memory[2445] = 12'h000;
    assign memory[2446] = 12'h000;
    assign memory[2447] = 12'h000;
    assign memory[2448] = 12'h000;
    assign memory[2449] = 12'h000;
    assign memory[2450] = 12'h000;
    assign memory[2451] = 12'h000;
    assign memory[2452] = 12'h000;
    assign memory[2453] = 12'h000;
    assign memory[2454] = 12'h000;
    assign memory[2455] = 12'h000;
    assign memory[2456] = 12'h000;
    assign memory[2457] = 12'h000;
    assign memory[2458] = 12'h000;
    assign memory[2459] = 12'h000;
    assign memory[2460] = 12'h000;
    assign memory[2461] = 12'h000;
    assign memory[2462] = 12'h000;
    assign memory[2463] = 12'h000;
    assign memory[2464] = 12'h000;
    assign memory[2465] = 12'h000;
    assign memory[2466] = 12'h000;
    assign memory[2467] = 12'h000;
    assign memory[2468] = 12'h000;
    assign memory[2469] = 12'h000;
    assign memory[2470] = 12'h000;
    assign memory[2471] = 12'h000;
    assign memory[2472] = 12'h000;
    assign memory[2473] = 12'h000;
    assign memory[2474] = 12'h000;
    assign memory[2475] = 12'h000;
    assign memory[2476] = 12'h000;
    assign memory[2477] = 12'h000;
    assign memory[2478] = 12'h000;
    assign memory[2479] = 12'h000;
    assign memory[2480] = 12'h000;
    assign memory[2481] = 12'h000;
    assign memory[2482] = 12'h000;
    assign memory[2483] = 12'h000;
    assign memory[2484] = 12'h000;
    assign memory[2485] = 12'h000;
    assign memory[2486] = 12'h000;
    assign memory[2487] = 12'h000;
    assign memory[2488] = 12'h000;
    assign memory[2489] = 12'h000;
    assign memory[2490] = 12'h000;
    assign memory[2491] = 12'h000;
    assign memory[2492] = 12'h000;
    assign memory[2493] = 12'h000;
    assign memory[2494] = 12'h000;
    assign memory[2495] = 12'h000;
    assign memory[2496] = 12'h000;
    assign memory[2497] = 12'h000;
    assign memory[2498] = 12'h000;
    assign memory[2499] = 12'h000;
    assign memory[2500] = 12'h000;
    assign memory[2501] = 12'h000;
    assign memory[2502] = 12'h000;
    assign memory[2503] = 12'h000;
    assign memory[2504] = 12'h000;
    assign memory[2505] = 12'h000;
    assign memory[2506] = 12'h000;
    assign memory[2507] = 12'h000;
    assign memory[2508] = 12'h000;
    assign memory[2509] = 12'h000;
    assign memory[2510] = 12'h000;
    assign memory[2511] = 12'h000;
    assign memory[2512] = 12'h000;
    assign memory[2513] = 12'h000;
    assign memory[2514] = 12'h000;
    assign memory[2515] = 12'h000;
    assign memory[2516] = 12'h000;
    assign memory[2517] = 12'h000;
    assign memory[2518] = 12'h000;
    assign memory[2519] = 12'h000;
    assign memory[2520] = 12'h000;
    assign memory[2521] = 12'h000;
    assign memory[2522] = 12'h000;
    assign memory[2523] = 12'h000;
    assign memory[2524] = 12'h000;
    assign memory[2525] = 12'h000;
    assign memory[2526] = 12'h000;
    assign memory[2527] = 12'h000;
    assign memory[2528] = 12'h000;
    assign memory[2529] = 12'h000;
    assign memory[2530] = 12'h000;
    assign memory[2531] = 12'h000;
    assign memory[2532] = 12'h000;
    assign memory[2533] = 12'h000;
    assign memory[2534] = 12'h000;
    assign memory[2535] = 12'h000;
    assign memory[2536] = 12'h000;
    assign memory[2537] = 12'h000;
    assign memory[2538] = 12'h000;
    assign memory[2539] = 12'h000;
    assign memory[2540] = 12'h000;
    assign memory[2541] = 12'h000;
    assign memory[2542] = 12'h000;
    assign memory[2543] = 12'h000;
    assign memory[2544] = 12'h000;
    assign memory[2545] = 12'h000;
    assign memory[2546] = 12'h000;
    assign memory[2547] = 12'h000;
    assign memory[2548] = 12'h000;
    assign memory[2549] = 12'h000;
    assign memory[2550] = 12'h000;
    assign memory[2551] = 12'h000;
    assign memory[2552] = 12'h000;
    assign memory[2553] = 12'h000;
    assign memory[2554] = 12'h000;
    assign memory[2555] = 12'h000;
    assign memory[2556] = 12'h000;
    assign memory[2557] = 12'h000;
    assign memory[2558] = 12'h000;
    assign memory[2559] = 12'h000;
    assign memory[2560] = 12'h000;
    assign memory[2561] = 12'h000;
    assign memory[2562] = 12'h000;
    assign memory[2563] = 12'h000;
    assign memory[2564] = 12'h000;
    assign memory[2565] = 12'h000;
    assign memory[2566] = 12'h000;
    assign memory[2567] = 12'h000;
    assign memory[2568] = 12'h000;
    assign memory[2569] = 12'h000;
    assign memory[2570] = 12'h000;
    assign memory[2571] = 12'h000;
    assign memory[2572] = 12'h000;
    assign memory[2573] = 12'h000;
    assign memory[2574] = 12'h000;
    assign memory[2575] = 12'h000;
    assign memory[2576] = 12'h000;
    assign memory[2577] = 12'h000;
    assign memory[2578] = 12'h000;
    assign memory[2579] = 12'h000;
    assign memory[2580] = 12'h000;
    assign memory[2581] = 12'h000;
    assign memory[2582] = 12'h000;
    assign memory[2583] = 12'h000;
    assign memory[2584] = 12'h000;
    assign memory[2585] = 12'h000;
    assign memory[2586] = 12'h000;
    assign memory[2587] = 12'h000;
    assign memory[2588] = 12'h000;
    assign memory[2589] = 12'h000;
    assign memory[2590] = 12'h000;
    assign memory[2591] = 12'h000;
    assign memory[2592] = 12'h000;
    assign memory[2593] = 12'h000;
    assign memory[2594] = 12'h000;
    assign memory[2595] = 12'h000;
    assign memory[2596] = 12'h000;
    assign memory[2597] = 12'h000;
    assign memory[2598] = 12'h000;
    assign memory[2599] = 12'h000;
    assign memory[2600] = 12'h000;
    assign memory[2601] = 12'h000;
    assign memory[2602] = 12'h000;
    assign memory[2603] = 12'h000;
    assign memory[2604] = 12'h000;
    assign memory[2605] = 12'h000;
    assign memory[2606] = 12'h000;
    assign memory[2607] = 12'h000;
    assign memory[2608] = 12'h000;
    assign memory[2609] = 12'h000;
    assign memory[2610] = 12'h000;
    assign memory[2611] = 12'h000;
    assign memory[2612] = 12'h000;
    assign memory[2613] = 12'h000;
    assign memory[2614] = 12'h000;
    assign memory[2615] = 12'h000;
    assign memory[2616] = 12'h000;
    assign memory[2617] = 12'h000;
    assign memory[2618] = 12'h000;
    assign memory[2619] = 12'h000;
    assign memory[2620] = 12'h000;
    assign memory[2621] = 12'h000;
    assign memory[2622] = 12'h000;
    assign memory[2623] = 12'h000;
    assign memory[2624] = 12'h000;
    assign memory[2625] = 12'h000;
    assign memory[2626] = 12'h000;
    assign memory[2627] = 12'h000;
    assign memory[2628] = 12'h000;
    assign memory[2629] = 12'h000;
    assign memory[2630] = 12'h000;
    assign memory[2631] = 12'h000;
    assign memory[2632] = 12'h000;
    assign memory[2633] = 12'h000;
    assign memory[2634] = 12'h000;
    assign memory[2635] = 12'h000;
    assign memory[2636] = 12'h000;
    assign memory[2637] = 12'h000;
    assign memory[2638] = 12'h000;
    assign memory[2639] = 12'h000;
    assign memory[2640] = 12'h000;
    assign memory[2641] = 12'h000;
    assign memory[2642] = 12'h000;
    assign memory[2643] = 12'h000;
    assign memory[2644] = 12'h000;
    assign memory[2645] = 12'h000;
    assign memory[2646] = 12'h000;
    assign memory[2647] = 12'h000;
    assign memory[2648] = 12'h000;
    assign memory[2649] = 12'h000;
    assign memory[2650] = 12'h000;
    assign memory[2651] = 12'h000;
    assign memory[2652] = 12'h000;
    assign memory[2653] = 12'h000;
    assign memory[2654] = 12'h000;
    assign memory[2655] = 12'h000;
    assign memory[2656] = 12'h000;
    assign memory[2657] = 12'h000;
    assign memory[2658] = 12'h000;
    assign memory[2659] = 12'h000;
    assign memory[2660] = 12'h000;
    assign memory[2661] = 12'h000;
    assign memory[2662] = 12'h000;
    assign memory[2663] = 12'h000;
    assign memory[2664] = 12'h000;
    assign memory[2665] = 12'h000;
    assign memory[2666] = 12'h000;
    assign memory[2667] = 12'h000;
    assign memory[2668] = 12'h000;
    assign memory[2669] = 12'h000;
    assign memory[2670] = 12'h000;
    assign memory[2671] = 12'h000;
    assign memory[2672] = 12'h000;
    assign memory[2673] = 12'h000;
    assign memory[2674] = 12'h000;
    assign memory[2675] = 12'h000;
    assign memory[2676] = 12'h000;
    assign memory[2677] = 12'h000;
    assign memory[2678] = 12'h000;
    assign memory[2679] = 12'h000;
    assign memory[2680] = 12'h000;
    assign memory[2681] = 12'h000;
    assign memory[2682] = 12'h000;
    assign memory[2683] = 12'h000;
    assign memory[2684] = 12'h000;
    assign memory[2685] = 12'h000;
    assign memory[2686] = 12'h000;
    assign memory[2687] = 12'h000;
    assign memory[2688] = 12'h000;
    assign memory[2689] = 12'h000;
    assign memory[2690] = 12'h000;
    assign memory[2691] = 12'h000;
    assign memory[2692] = 12'h000;
    assign memory[2693] = 12'h000;
    assign memory[2694] = 12'h000;
    assign memory[2695] = 12'h000;
    assign memory[2696] = 12'h000;
    assign memory[2697] = 12'h000;
    assign memory[2698] = 12'h000;
    assign memory[2699] = 12'h000;
    assign memory[2700] = 12'h000;
    assign memory[2701] = 12'h000;
    assign memory[2702] = 12'h000;
    assign memory[2703] = 12'h000;
    assign memory[2704] = 12'h000;
    assign memory[2705] = 12'h000;
    assign memory[2706] = 12'h000;
    assign memory[2707] = 12'h000;
    assign memory[2708] = 12'h000;
    assign memory[2709] = 12'h000;
    assign memory[2710] = 12'h000;
    assign memory[2711] = 12'h000;
    assign memory[2712] = 12'h000;
    assign memory[2713] = 12'h000;
    assign memory[2714] = 12'h000;
    assign memory[2715] = 12'h000;
    assign memory[2716] = 12'h000;
    assign memory[2717] = 12'h000;
    assign memory[2718] = 12'h000;
    assign memory[2719] = 12'h000;
    assign memory[2720] = 12'h000;
    assign memory[2721] = 12'h000;
    assign memory[2722] = 12'h000;
    assign memory[2723] = 12'h000;
    assign memory[2724] = 12'h000;
    assign memory[2725] = 12'h000;
    assign memory[2726] = 12'h000;
    assign memory[2727] = 12'h000;
    assign memory[2728] = 12'h000;
    assign memory[2729] = 12'h000;
    assign memory[2730] = 12'h000;
    assign memory[2731] = 12'h000;
    assign memory[2732] = 12'h000;
    assign memory[2733] = 12'h000;
    assign memory[2734] = 12'h000;
    assign memory[2735] = 12'h000;
    assign memory[2736] = 12'h000;
    assign memory[2737] = 12'h000;
    assign memory[2738] = 12'h000;
    assign memory[2739] = 12'h000;
    assign memory[2740] = 12'h000;
    assign memory[2741] = 12'h000;
    assign memory[2742] = 12'h000;
    assign memory[2743] = 12'h000;
    assign memory[2744] = 12'h000;
    assign memory[2745] = 12'h000;
    assign memory[2746] = 12'h000;
    assign memory[2747] = 12'h000;
    assign memory[2748] = 12'h000;
    assign memory[2749] = 12'h000;
    assign memory[2750] = 12'h000;
    assign memory[2751] = 12'h000;
    assign memory[2752] = 12'h000;
    assign memory[2753] = 12'h000;
    assign memory[2754] = 12'h000;
    assign memory[2755] = 12'h000;
    assign memory[2756] = 12'h000;
    assign memory[2757] = 12'h000;
    assign memory[2758] = 12'h000;
    assign memory[2759] = 12'h000;
    assign memory[2760] = 12'h000;
    assign memory[2761] = 12'h000;
    assign memory[2762] = 12'h000;
    assign memory[2763] = 12'h000;
    assign memory[2764] = 12'h000;
    assign memory[2765] = 12'h000;
    assign memory[2766] = 12'h000;
    assign memory[2767] = 12'h000;
    assign memory[2768] = 12'h000;
    assign memory[2769] = 12'h000;
    assign memory[2770] = 12'h000;
    assign memory[2771] = 12'h000;
    assign memory[2772] = 12'h000;
    assign memory[2773] = 12'h000;
    assign memory[2774] = 12'h000;
    assign memory[2775] = 12'h000;
    assign memory[2776] = 12'h000;
    assign memory[2777] = 12'h000;
    assign memory[2778] = 12'h000;
    assign memory[2779] = 12'h000;
    assign memory[2780] = 12'h000;
    assign memory[2781] = 12'h000;
    assign memory[2782] = 12'h000;
    assign memory[2783] = 12'h000;
    assign memory[2784] = 12'h000;
    assign memory[2785] = 12'h000;
    assign memory[2786] = 12'h000;
    assign memory[2787] = 12'h000;
    assign memory[2788] = 12'h000;
    assign memory[2789] = 12'h000;
    assign memory[2790] = 12'h000;
    assign memory[2791] = 12'h000;
    assign memory[2792] = 12'h000;
    assign memory[2793] = 12'h000;
    assign memory[2794] = 12'h000;
    assign memory[2795] = 12'h000;
    assign memory[2796] = 12'h000;
    assign memory[2797] = 12'h000;
    assign memory[2798] = 12'h000;
    assign memory[2799] = 12'h000;
    assign memory[2800] = 12'h000;
    assign memory[2801] = 12'h000;
    assign memory[2802] = 12'h000;
    assign memory[2803] = 12'h000;
    assign memory[2804] = 12'h000;
    assign memory[2805] = 12'h000;
    assign memory[2806] = 12'h000;
    assign memory[2807] = 12'h000;
    assign memory[2808] = 12'h000;
    assign memory[2809] = 12'h000;
    assign memory[2810] = 12'h000;
    assign memory[2811] = 12'h000;
    assign memory[2812] = 12'h000;
    assign memory[2813] = 12'h000;
    assign memory[2814] = 12'h000;
    assign memory[2815] = 12'h000;
    assign memory[2816] = 12'h000;
    assign memory[2817] = 12'h000;
    assign memory[2818] = 12'h000;
    assign memory[2819] = 12'h000;
    assign memory[2820] = 12'h000;
    assign memory[2821] = 12'h000;
    assign memory[2822] = 12'h000;
    assign memory[2823] = 12'h000;
    assign memory[2824] = 12'h000;
    assign memory[2825] = 12'h000;
    assign memory[2826] = 12'h000;
    assign memory[2827] = 12'h000;
    assign memory[2828] = 12'h000;
    assign memory[2829] = 12'h000;
    assign memory[2830] = 12'h000;
    assign memory[2831] = 12'h000;
    assign memory[2832] = 12'h000;
    assign memory[2833] = 12'h000;
    assign memory[2834] = 12'h000;
    assign memory[2835] = 12'h000;
    assign memory[2836] = 12'h000;
    assign memory[2837] = 12'h000;
    assign memory[2838] = 12'h000;
    assign memory[2839] = 12'h000;
    assign memory[2840] = 12'h000;
    assign memory[2841] = 12'h000;
    assign memory[2842] = 12'h000;
    assign memory[2843] = 12'h000;
    assign memory[2844] = 12'h000;
    assign memory[2845] = 12'h000;
    assign memory[2846] = 12'h000;
    assign memory[2847] = 12'h000;
    assign memory[2848] = 12'h000;
    assign memory[2849] = 12'h000;
    assign memory[2850] = 12'h000;
    assign memory[2851] = 12'h000;
    assign memory[2852] = 12'h000;
    assign memory[2853] = 12'h000;
    assign memory[2854] = 12'h000;
    assign memory[2855] = 12'h000;
    assign memory[2856] = 12'h000;
    assign memory[2857] = 12'h000;
    assign memory[2858] = 12'h000;
    assign memory[2859] = 12'h000;
    assign memory[2860] = 12'h000;
    assign memory[2861] = 12'h000;
    assign memory[2862] = 12'h000;
    assign memory[2863] = 12'h000;
    assign memory[2864] = 12'h000;
    assign memory[2865] = 12'h000;
    assign memory[2866] = 12'h000;
    assign memory[2867] = 12'h000;
    assign memory[2868] = 12'h000;
    assign memory[2869] = 12'h000;
    assign memory[2870] = 12'h000;
    assign memory[2871] = 12'h000;
    assign memory[2872] = 12'h000;
    assign memory[2873] = 12'h000;
    assign memory[2874] = 12'h000;
    assign memory[2875] = 12'h000;
    assign memory[2876] = 12'h000;
    assign memory[2877] = 12'h000;
    assign memory[2878] = 12'h000;
    assign memory[2879] = 12'h000;
    assign memory[2880] = 12'h000;
    assign memory[2881] = 12'h000;
    assign memory[2882] = 12'h000;
    assign memory[2883] = 12'h000;
    assign memory[2884] = 12'h000;
    assign memory[2885] = 12'h000;
    assign memory[2886] = 12'h000;
    assign memory[2887] = 12'h000;
    assign memory[2888] = 12'h000;
    assign memory[2889] = 12'h000;
    assign memory[2890] = 12'h000;
    assign memory[2891] = 12'h000;
    assign memory[2892] = 12'h000;
    assign memory[2893] = 12'h000;
    assign memory[2894] = 12'h000;
    assign memory[2895] = 12'h000;
    assign memory[2896] = 12'h000;
    assign memory[2897] = 12'h000;
    assign memory[2898] = 12'h000;
    assign memory[2899] = 12'h000;
    assign memory[2900] = 12'h000;
    assign memory[2901] = 12'h000;
    assign memory[2902] = 12'h000;
    assign memory[2903] = 12'h000;
    assign memory[2904] = 12'h000;
    assign memory[2905] = 12'h000;
    assign memory[2906] = 12'h000;
    assign memory[2907] = 12'h000;
    assign memory[2908] = 12'h000;
    assign memory[2909] = 12'h000;
    assign memory[2910] = 12'h000;
    assign memory[2911] = 12'h000;
    assign memory[2912] = 12'h000;
    assign memory[2913] = 12'h000;
    assign memory[2914] = 12'h000;
    assign memory[2915] = 12'h000;
    assign memory[2916] = 12'h000;
    assign memory[2917] = 12'h000;
    assign memory[2918] = 12'h000;
    assign memory[2919] = 12'h000;
    assign memory[2920] = 12'h000;
    assign memory[2921] = 12'h000;
    assign memory[2922] = 12'h000;
    assign memory[2923] = 12'h000;
    assign memory[2924] = 12'h000;
    assign memory[2925] = 12'h000;
    assign memory[2926] = 12'h000;
    assign memory[2927] = 12'h000;
    assign memory[2928] = 12'h000;
    assign memory[2929] = 12'h000;
    assign memory[2930] = 12'h000;
    assign memory[2931] = 12'h000;
    assign memory[2932] = 12'h000;
    assign memory[2933] = 12'h000;
    assign memory[2934] = 12'h000;
    assign memory[2935] = 12'h000;
    assign memory[2936] = 12'h000;
    assign memory[2937] = 12'h000;
    assign memory[2938] = 12'h000;
    assign memory[2939] = 12'h000;
    assign memory[2940] = 12'h000;
    assign memory[2941] = 12'h000;
    assign memory[2942] = 12'h000;
    assign memory[2943] = 12'h000;
    assign memory[2944] = 12'h000;
    assign memory[2945] = 12'h000;
    assign memory[2946] = 12'h000;
    assign memory[2947] = 12'h000;
    assign memory[2948] = 12'h000;
    assign memory[2949] = 12'h000;
    assign memory[2950] = 12'h000;
    assign memory[2951] = 12'h000;
    assign memory[2952] = 12'h000;
    assign memory[2953] = 12'h000;
    assign memory[2954] = 12'h000;
    assign memory[2955] = 12'h000;
    assign memory[2956] = 12'h000;
    assign memory[2957] = 12'h000;
    assign memory[2958] = 12'h000;
    assign memory[2959] = 12'h000;
    assign memory[2960] = 12'h000;
    assign memory[2961] = 12'h000;
    assign memory[2962] = 12'h000;
    assign memory[2963] = 12'h000;
    assign memory[2964] = 12'h000;
    assign memory[2965] = 12'h000;
    assign memory[2966] = 12'h000;
    assign memory[2967] = 12'h000;
    assign memory[2968] = 12'h000;
    assign memory[2969] = 12'h000;
    assign memory[2970] = 12'h000;
    assign memory[2971] = 12'h000;
    assign memory[2972] = 12'h000;
    assign memory[2973] = 12'h000;
    assign memory[2974] = 12'h000;
    assign memory[2975] = 12'h000;
    assign memory[2976] = 12'h000;
    assign memory[2977] = 12'h000;
    assign memory[2978] = 12'h000;
    assign memory[2979] = 12'h000;
    assign memory[2980] = 12'h000;
    assign memory[2981] = 12'h000;
    assign memory[2982] = 12'h000;
    assign memory[2983] = 12'h000;
    assign memory[2984] = 12'h000;
    assign memory[2985] = 12'h000;
    assign memory[2986] = 12'h000;
    assign memory[2987] = 12'h000;
    assign memory[2988] = 12'h000;
    assign memory[2989] = 12'h000;
    assign memory[2990] = 12'h000;
    assign memory[2991] = 12'h000;
    assign memory[2992] = 12'h000;
    assign memory[2993] = 12'h000;
    assign memory[2994] = 12'h000;
    assign memory[2995] = 12'h000;
    assign memory[2996] = 12'h000;
    assign memory[2997] = 12'h000;
    assign memory[2998] = 12'h000;
    assign memory[2999] = 12'h000;
    assign memory[3000] = 12'h000;
    assign memory[3001] = 12'h000;
    assign memory[3002] = 12'h000;
    assign memory[3003] = 12'h000;
    assign memory[3004] = 12'h000;
    assign memory[3005] = 12'h000;
    assign memory[3006] = 12'h000;
    assign memory[3007] = 12'h000;
    assign memory[3008] = 12'h000;
    assign memory[3009] = 12'h000;
    assign memory[3010] = 12'h000;
    assign memory[3011] = 12'h000;
    assign memory[3012] = 12'h000;
    assign memory[3013] = 12'h000;
    assign memory[3014] = 12'h000;
    assign memory[3015] = 12'h000;
    assign memory[3016] = 12'h000;
    assign memory[3017] = 12'h000;
    assign memory[3018] = 12'h000;
    assign memory[3019] = 12'h000;
    assign memory[3020] = 12'h000;
    assign memory[3021] = 12'h000;
    assign memory[3022] = 12'h000;
    assign memory[3023] = 12'h000;
    assign memory[3024] = 12'h000;
    assign memory[3025] = 12'h000;
    assign memory[3026] = 12'h000;
    assign memory[3027] = 12'h000;
    assign memory[3028] = 12'h000;
    assign memory[3029] = 12'h000;
    assign memory[3030] = 12'h000;
    assign memory[3031] = 12'h000;
    assign memory[3032] = 12'h000;
    assign memory[3033] = 12'h000;
    assign memory[3034] = 12'h000;
    assign memory[3035] = 12'h000;
    assign memory[3036] = 12'h000;
    assign memory[3037] = 12'h000;
    assign memory[3038] = 12'h000;
    assign memory[3039] = 12'h000;
    assign memory[3040] = 12'h000;
    assign memory[3041] = 12'h000;
    assign memory[3042] = 12'h000;
    assign memory[3043] = 12'h000;
    assign memory[3044] = 12'h000;
    assign memory[3045] = 12'h000;
    assign memory[3046] = 12'h000;
    assign memory[3047] = 12'h000;
    assign memory[3048] = 12'h000;
    assign memory[3049] = 12'h000;
    assign memory[3050] = 12'h000;
    assign memory[3051] = 12'h000;
    assign memory[3052] = 12'h000;
    assign memory[3053] = 12'h000;
    assign memory[3054] = 12'h000;
    assign memory[3055] = 12'h000;
    assign memory[3056] = 12'h000;
    assign memory[3057] = 12'h000;
    assign memory[3058] = 12'h000;
    assign memory[3059] = 12'h000;
    assign memory[3060] = 12'h000;
    assign memory[3061] = 12'h000;
    assign memory[3062] = 12'h000;
    assign memory[3063] = 12'h000;
    assign memory[3064] = 12'h000;
    assign memory[3065] = 12'h000;
    assign memory[3066] = 12'h000;
    assign memory[3067] = 12'h000;
    assign memory[3068] = 12'h000;
    assign memory[3069] = 12'h000;
    assign memory[3070] = 12'h000;
    assign memory[3071] = 12'h000;
    assign memory[3072] = 12'hfff;
    assign memory[3073] = 12'hfff;
    assign memory[3074] = 12'hfff;
    assign memory[3075] = 12'hfff;
    assign memory[3076] = 12'hfff;
    assign memory[3077] = 12'hfff;
    assign memory[3078] = 12'hfff;
    assign memory[3079] = 12'hfff;
    assign memory[3080] = 12'hfff;
    assign memory[3081] = 12'hfff;
    assign memory[3082] = 12'hfff;
    assign memory[3083] = 12'hfff;
    assign memory[3084] = 12'hfff;
    assign memory[3085] = 12'hfff;
    assign memory[3086] = 12'hfff;
    assign memory[3087] = 12'hfff;
    assign memory[3088] = 12'hfff;
    assign memory[3089] = 12'hfff;
    assign memory[3090] = 12'hfff;
    assign memory[3091] = 12'hfff;
    assign memory[3092] = 12'hfff;
    assign memory[3093] = 12'hfff;
    assign memory[3094] = 12'hfff;
    assign memory[3095] = 12'hfff;
    assign memory[3096] = 12'hfff;
    assign memory[3097] = 12'hfff;
    assign memory[3098] = 12'hfff;
    assign memory[3099] = 12'hfff;
    assign memory[3100] = 12'hfff;
    assign memory[3101] = 12'hfff;
    assign memory[3102] = 12'hfff;
    assign memory[3103] = 12'hfff;
    assign memory[3104] = 12'hfff;
    assign memory[3105] = 12'hfff;
    assign memory[3106] = 12'hfff;
    assign memory[3107] = 12'hfff;
    assign memory[3108] = 12'hfff;
    assign memory[3109] = 12'hfff;
    assign memory[3110] = 12'hfff;
    assign memory[3111] = 12'hfff;
    assign memory[3112] = 12'hfff;
    assign memory[3113] = 12'hfff;
    assign memory[3114] = 12'hfff;
    assign memory[3115] = 12'hfff;
    assign memory[3116] = 12'hfff;
    assign memory[3117] = 12'hfff;
    assign memory[3118] = 12'hfff;
    assign memory[3119] = 12'hfff;
    assign memory[3120] = 12'hfff;
    assign memory[3121] = 12'hfff;
    assign memory[3122] = 12'hfff;
    assign memory[3123] = 12'hfff;
    assign memory[3124] = 12'hfff;
    assign memory[3125] = 12'hfff;
    assign memory[3126] = 12'hfff;
    assign memory[3127] = 12'hfff;
    assign memory[3128] = 12'hfff;
    assign memory[3129] = 12'hfff;
    assign memory[3130] = 12'hfff;
    assign memory[3131] = 12'hfff;
    assign memory[3132] = 12'hfff;
    assign memory[3133] = 12'hfff;
    assign memory[3134] = 12'hfff;
    assign memory[3135] = 12'hfff;
    assign memory[3136] = 12'hfff;
    assign memory[3137] = 12'hfff;
    assign memory[3138] = 12'hfff;
    assign memory[3139] = 12'hfff;
    assign memory[3140] = 12'hfff;
    assign memory[3141] = 12'hfff;
    assign memory[3142] = 12'hfff;
    assign memory[3143] = 12'hfff;
    assign memory[3144] = 12'hfff;
    assign memory[3145] = 12'hfff;
    assign memory[3146] = 12'hfff;
    assign memory[3147] = 12'hfff;
    assign memory[3148] = 12'hfff;
    assign memory[3149] = 12'hfff;
    assign memory[3150] = 12'hfff;
    assign memory[3151] = 12'hfff;
    assign memory[3152] = 12'hfff;
    assign memory[3153] = 12'hfff;
    assign memory[3154] = 12'hfff;
    assign memory[3155] = 12'hfff;
    assign memory[3156] = 12'hfff;
    assign memory[3157] = 12'hfff;
    assign memory[3158] = 12'hfff;
    assign memory[3159] = 12'hfff;
    assign memory[3160] = 12'hfff;
    assign memory[3161] = 12'hfff;
    assign memory[3162] = 12'hfff;
    assign memory[3163] = 12'hfff;
    assign memory[3164] = 12'hfff;
    assign memory[3165] = 12'hfff;
    assign memory[3166] = 12'hfff;
    assign memory[3167] = 12'hfff;
    assign memory[3168] = 12'hfff;
    assign memory[3169] = 12'hfff;
    assign memory[3170] = 12'hfff;
    assign memory[3171] = 12'hfff;
    assign memory[3172] = 12'hfff;
    assign memory[3173] = 12'hfff;
    assign memory[3174] = 12'hfff;
    assign memory[3175] = 12'hfff;
    assign memory[3176] = 12'hfff;
    assign memory[3177] = 12'hfff;
    assign memory[3178] = 12'hfff;
    assign memory[3179] = 12'hfff;
    assign memory[3180] = 12'hfff;
    assign memory[3181] = 12'hfff;
    assign memory[3182] = 12'hfff;
    assign memory[3183] = 12'hfff;
    assign memory[3184] = 12'hfff;
    assign memory[3185] = 12'hfff;
    assign memory[3186] = 12'hfff;
    assign memory[3187] = 12'hfff;
    assign memory[3188] = 12'hfff;
    assign memory[3189] = 12'hfff;
    assign memory[3190] = 12'hfff;
    assign memory[3191] = 12'hfff;
    assign memory[3192] = 12'hfff;
    assign memory[3193] = 12'hfff;
    assign memory[3194] = 12'hfff;
    assign memory[3195] = 12'hfff;
    assign memory[3196] = 12'hfff;
    assign memory[3197] = 12'hfff;
    assign memory[3198] = 12'hfff;
    assign memory[3199] = 12'hfff;
    assign memory[3200] = 12'hfff;
    assign memory[3201] = 12'hfff;
    assign memory[3202] = 12'hfff;
    assign memory[3203] = 12'hfff;
    assign memory[3204] = 12'hfff;
    assign memory[3205] = 12'hfff;
    assign memory[3206] = 12'hfff;
    assign memory[3207] = 12'hfff;
    assign memory[3208] = 12'hfff;
    assign memory[3209] = 12'hfff;
    assign memory[3210] = 12'hfff;
    assign memory[3211] = 12'hfff;
    assign memory[3212] = 12'hfff;
    assign memory[3213] = 12'hfff;
    assign memory[3214] = 12'hfff;
    assign memory[3215] = 12'hfff;
    assign memory[3216] = 12'hfff;
    assign memory[3217] = 12'hfff;
    assign memory[3218] = 12'hfff;
    assign memory[3219] = 12'hfff;
    assign memory[3220] = 12'hfff;
    assign memory[3221] = 12'hfff;
    assign memory[3222] = 12'hfff;
    assign memory[3223] = 12'hfff;
    assign memory[3224] = 12'hfff;
    assign memory[3225] = 12'hfff;
    assign memory[3226] = 12'hfff;
    assign memory[3227] = 12'hfff;
    assign memory[3228] = 12'hfff;
    assign memory[3229] = 12'hfff;
    assign memory[3230] = 12'hfff;
    assign memory[3231] = 12'hfff;
    assign memory[3232] = 12'hfff;
    assign memory[3233] = 12'hfff;
    assign memory[3234] = 12'hfff;
    assign memory[3235] = 12'hfff;
    assign memory[3236] = 12'hfff;
    assign memory[3237] = 12'hfff;
    assign memory[3238] = 12'hfff;
    assign memory[3239] = 12'hfff;
    assign memory[3240] = 12'hfff;
    assign memory[3241] = 12'hfff;
    assign memory[3242] = 12'hfff;
    assign memory[3243] = 12'hfff;
    assign memory[3244] = 12'hfff;
    assign memory[3245] = 12'hfff;
    assign memory[3246] = 12'hfff;
    assign memory[3247] = 12'hfff;
    assign memory[3248] = 12'hfff;
    assign memory[3249] = 12'hfff;
    assign memory[3250] = 12'hfff;
    assign memory[3251] = 12'hfff;
    assign memory[3252] = 12'hfff;
    assign memory[3253] = 12'hfff;
    assign memory[3254] = 12'hfff;
    assign memory[3255] = 12'hfff;
    assign memory[3256] = 12'hfff;
    assign memory[3257] = 12'hfff;
    assign memory[3258] = 12'hfff;
    assign memory[3259] = 12'hfff;
    assign memory[3260] = 12'hfff;
    assign memory[3261] = 12'hfff;
    assign memory[3262] = 12'hfff;
    assign memory[3263] = 12'hfff;
    assign memory[3264] = 12'hfff;
    assign memory[3265] = 12'hfff;
    assign memory[3266] = 12'hfff;
    assign memory[3267] = 12'hfff;
    assign memory[3268] = 12'hfff;
    assign memory[3269] = 12'hfff;
    assign memory[3270] = 12'hfff;
    assign memory[3271] = 12'hfff;
    assign memory[3272] = 12'hfff;
    assign memory[3273] = 12'hfff;
    assign memory[3274] = 12'hfff;
    assign memory[3275] = 12'hfff;
    assign memory[3276] = 12'hfff;
    assign memory[3277] = 12'hfff;
    assign memory[3278] = 12'hfff;
    assign memory[3279] = 12'hfff;
    assign memory[3280] = 12'hfff;
    assign memory[3281] = 12'hfff;
    assign memory[3282] = 12'hfff;
    assign memory[3283] = 12'hfff;
    assign memory[3284] = 12'hfff;
    assign memory[3285] = 12'hfff;
    assign memory[3286] = 12'hfff;
    assign memory[3287] = 12'hfff;
    assign memory[3288] = 12'hfff;
    assign memory[3289] = 12'hfff;
    assign memory[3290] = 12'hfff;
    assign memory[3291] = 12'hfff;
    assign memory[3292] = 12'hfff;
    assign memory[3293] = 12'hfff;
    assign memory[3294] = 12'hfff;
    assign memory[3295] = 12'hfff;
    assign memory[3296] = 12'hfff;
    assign memory[3297] = 12'hfff;
    assign memory[3298] = 12'hfff;
    assign memory[3299] = 12'hfff;
    assign memory[3300] = 12'hfff;
    assign memory[3301] = 12'hfff;
    assign memory[3302] = 12'hfff;
    assign memory[3303] = 12'hfff;
    assign memory[3304] = 12'hfff;
    assign memory[3305] = 12'hfff;
    assign memory[3306] = 12'hfff;
    assign memory[3307] = 12'hfff;
    assign memory[3308] = 12'hfff;
    assign memory[3309] = 12'hfff;
    assign memory[3310] = 12'hfff;
    assign memory[3311] = 12'hfff;
    assign memory[3312] = 12'hfff;
    assign memory[3313] = 12'hfff;
    assign memory[3314] = 12'hfff;
    assign memory[3315] = 12'hfff;
    assign memory[3316] = 12'hfff;
    assign memory[3317] = 12'hfff;
    assign memory[3318] = 12'hfff;
    assign memory[3319] = 12'hfff;
    assign memory[3320] = 12'hfff;
    assign memory[3321] = 12'hfff;
    assign memory[3322] = 12'hfff;
    assign memory[3323] = 12'hfff;
    assign memory[3324] = 12'hfff;
    assign memory[3325] = 12'hfff;
    assign memory[3326] = 12'hfff;
    assign memory[3327] = 12'hfff;
    assign memory[3328] = 12'hfff;
    assign memory[3329] = 12'hfff;
    assign memory[3330] = 12'hfff;
    assign memory[3331] = 12'hfff;
    assign memory[3332] = 12'hfff;
    assign memory[3333] = 12'hfff;
    assign memory[3334] = 12'hfff;
    assign memory[3335] = 12'hfff;
    assign memory[3336] = 12'hfff;
    assign memory[3337] = 12'hfff;
    assign memory[3338] = 12'hfff;
    assign memory[3339] = 12'hfff;
    assign memory[3340] = 12'hfff;
    assign memory[3341] = 12'hfff;
    assign memory[3342] = 12'hfff;
    assign memory[3343] = 12'hfff;
    assign memory[3344] = 12'hfff;
    assign memory[3345] = 12'hfff;
    assign memory[3346] = 12'hfff;
    assign memory[3347] = 12'hfff;
    assign memory[3348] = 12'hfff;
    assign memory[3349] = 12'hfff;
    assign memory[3350] = 12'hfff;
    assign memory[3351] = 12'hfff;
    assign memory[3352] = 12'hfff;
    assign memory[3353] = 12'hfff;
    assign memory[3354] = 12'hfff;
    assign memory[3355] = 12'hfff;
    assign memory[3356] = 12'hfff;
    assign memory[3357] = 12'hfff;
    assign memory[3358] = 12'hfff;
    assign memory[3359] = 12'hfff;
    assign memory[3360] = 12'hfff;
    assign memory[3361] = 12'hfff;
    assign memory[3362] = 12'hfff;
    assign memory[3363] = 12'hfff;
    assign memory[3364] = 12'hfff;
    assign memory[3365] = 12'hfff;
    assign memory[3366] = 12'hfff;
    assign memory[3367] = 12'hfff;
    assign memory[3368] = 12'hfff;
    assign memory[3369] = 12'hfff;
    assign memory[3370] = 12'hfff;
    assign memory[3371] = 12'hfff;
    assign memory[3372] = 12'hfff;
    assign memory[3373] = 12'hfff;
    assign memory[3374] = 12'hfff;
    assign memory[3375] = 12'hfff;
    assign memory[3376] = 12'hfff;
    assign memory[3377] = 12'hfff;
    assign memory[3378] = 12'hfff;
    assign memory[3379] = 12'hfff;
    assign memory[3380] = 12'hfff;
    assign memory[3381] = 12'hfff;
    assign memory[3382] = 12'hfff;
    assign memory[3383] = 12'hfff;
    assign memory[3384] = 12'hfff;
    assign memory[3385] = 12'hfff;
    assign memory[3386] = 12'hfff;
    assign memory[3387] = 12'hfff;
    assign memory[3388] = 12'hfff;
    assign memory[3389] = 12'hfff;
    assign memory[3390] = 12'hfff;
    assign memory[3391] = 12'hfff;
    assign memory[3392] = 12'hfff;
    assign memory[3393] = 12'hfff;
    assign memory[3394] = 12'hfff;
    assign memory[3395] = 12'hfff;
    assign memory[3396] = 12'hfff;
    assign memory[3397] = 12'hfff;
    assign memory[3398] = 12'hfff;
    assign memory[3399] = 12'hfff;
    assign memory[3400] = 12'hfff;
    assign memory[3401] = 12'hfff;
    assign memory[3402] = 12'hfff;
    assign memory[3403] = 12'hfff;
    assign memory[3404] = 12'hfff;
    assign memory[3405] = 12'hfff;
    assign memory[3406] = 12'hfff;
    assign memory[3407] = 12'hfff;
    assign memory[3408] = 12'hfff;
    assign memory[3409] = 12'hfff;
    assign memory[3410] = 12'hfff;
    assign memory[3411] = 12'hfff;
    assign memory[3412] = 12'hfff;
    assign memory[3413] = 12'hfff;
    assign memory[3414] = 12'hfff;
    assign memory[3415] = 12'hfff;
    assign memory[3416] = 12'hfff;
    assign memory[3417] = 12'hfff;
    assign memory[3418] = 12'hfff;
    assign memory[3419] = 12'hfff;
    assign memory[3420] = 12'hfff;
    assign memory[3421] = 12'hfff;
    assign memory[3422] = 12'hfff;
    assign memory[3423] = 12'hfff;
    assign memory[3424] = 12'hfff;
    assign memory[3425] = 12'hfff;
    assign memory[3426] = 12'hfff;
    assign memory[3427] = 12'hfff;
    assign memory[3428] = 12'hfff;
    assign memory[3429] = 12'hfff;
    assign memory[3430] = 12'hfff;
    assign memory[3431] = 12'hfff;
    assign memory[3432] = 12'hfff;
    assign memory[3433] = 12'hfff;
    assign memory[3434] = 12'hfff;
    assign memory[3435] = 12'hfff;
    assign memory[3436] = 12'hfff;
    assign memory[3437] = 12'hfff;
    assign memory[3438] = 12'hfff;
    assign memory[3439] = 12'hfff;
    assign memory[3440] = 12'hfff;
    assign memory[3441] = 12'hfff;
    assign memory[3442] = 12'hfff;
    assign memory[3443] = 12'hfff;
    assign memory[3444] = 12'hfff;
    assign memory[3445] = 12'hfff;
    assign memory[3446] = 12'hfff;
    assign memory[3447] = 12'hfff;
    assign memory[3448] = 12'hfff;
    assign memory[3449] = 12'hfff;
    assign memory[3450] = 12'hfff;
    assign memory[3451] = 12'hfff;
    assign memory[3452] = 12'hfff;
    assign memory[3453] = 12'hfff;
    assign memory[3454] = 12'hfff;
    assign memory[3455] = 12'hfff;
    assign memory[3456] = 12'hfff;
    assign memory[3457] = 12'hfff;
    assign memory[3458] = 12'hfff;
    assign memory[3459] = 12'hfff;
    assign memory[3460] = 12'hfff;
    assign memory[3461] = 12'hfff;
    assign memory[3462] = 12'hfff;
    assign memory[3463] = 12'hfff;
    assign memory[3464] = 12'hfff;
    assign memory[3465] = 12'hfff;
    assign memory[3466] = 12'hfff;
    assign memory[3467] = 12'hfff;
    assign memory[3468] = 12'hfff;
    assign memory[3469] = 12'hfff;
    assign memory[3470] = 12'hfff;
    assign memory[3471] = 12'hfff;
    assign memory[3472] = 12'hfff;
    assign memory[3473] = 12'hfff;
    assign memory[3474] = 12'hfff;
    assign memory[3475] = 12'hfff;
    assign memory[3476] = 12'hfff;
    assign memory[3477] = 12'hfff;
    assign memory[3478] = 12'hfff;
    assign memory[3479] = 12'hfff;
    assign memory[3480] = 12'hfff;
    assign memory[3481] = 12'hfff;
    assign memory[3482] = 12'hfff;
    assign memory[3483] = 12'hfff;
    assign memory[3484] = 12'hfff;
    assign memory[3485] = 12'hfff;
    assign memory[3486] = 12'hfff;
    assign memory[3487] = 12'hfff;
    assign memory[3488] = 12'hfff;
    assign memory[3489] = 12'hfff;
    assign memory[3490] = 12'hfff;
    assign memory[3491] = 12'hfff;
    assign memory[3492] = 12'hfff;
    assign memory[3493] = 12'hfff;
    assign memory[3494] = 12'hfff;
    assign memory[3495] = 12'hfff;
    assign memory[3496] = 12'hfff;
    assign memory[3497] = 12'hfff;
    assign memory[3498] = 12'hfff;
    assign memory[3499] = 12'hfff;
    assign memory[3500] = 12'hfff;
    assign memory[3501] = 12'hfff;
    assign memory[3502] = 12'hfff;
    assign memory[3503] = 12'hfff;
    assign memory[3504] = 12'hfff;
    assign memory[3505] = 12'hfff;
    assign memory[3506] = 12'hfff;
    assign memory[3507] = 12'hfff;
    assign memory[3508] = 12'hfff;
    assign memory[3509] = 12'hfff;
    assign memory[3510] = 12'hfff;
    assign memory[3511] = 12'hfff;
    assign memory[3512] = 12'hfff;
    assign memory[3513] = 12'hfff;
    assign memory[3514] = 12'hfff;
    assign memory[3515] = 12'hfff;
    assign memory[3516] = 12'hfff;
    assign memory[3517] = 12'hfff;
    assign memory[3518] = 12'hfff;
    assign memory[3519] = 12'hfff;
    assign memory[3520] = 12'hfff;
    assign memory[3521] = 12'hfff;
    assign memory[3522] = 12'hfff;
    assign memory[3523] = 12'hfff;
    assign memory[3524] = 12'hfff;
    assign memory[3525] = 12'hfff;
    assign memory[3526] = 12'hfff;
    assign memory[3527] = 12'hfff;
    assign memory[3528] = 12'hfff;
    assign memory[3529] = 12'hfff;
    assign memory[3530] = 12'hfff;
    assign memory[3531] = 12'hfff;
    assign memory[3532] = 12'hfff;
    assign memory[3533] = 12'hfff;
    assign memory[3534] = 12'hfff;
    assign memory[3535] = 12'hfff;
    assign memory[3536] = 12'hfff;
    assign memory[3537] = 12'hfff;
    assign memory[3538] = 12'hfff;
    assign memory[3539] = 12'hfff;
    assign memory[3540] = 12'hfff;
    assign memory[3541] = 12'hfff;
    assign memory[3542] = 12'hfff;
    assign memory[3543] = 12'hfff;
    assign memory[3544] = 12'hfff;
    assign memory[3545] = 12'hfff;
    assign memory[3546] = 12'hfff;
    assign memory[3547] = 12'hfff;
    assign memory[3548] = 12'hfff;
    assign memory[3549] = 12'hfff;
    assign memory[3550] = 12'hfff;
    assign memory[3551] = 12'hfff;
    assign memory[3552] = 12'hfff;
    assign memory[3553] = 12'hfff;
    assign memory[3554] = 12'hfff;
    assign memory[3555] = 12'hfff;
    assign memory[3556] = 12'hfff;
    assign memory[3557] = 12'hfff;
    assign memory[3558] = 12'hfff;
    assign memory[3559] = 12'hfff;
    assign memory[3560] = 12'hfff;
    assign memory[3561] = 12'hfff;
    assign memory[3562] = 12'hfff;
    assign memory[3563] = 12'hfff;
    assign memory[3564] = 12'hfff;
    assign memory[3565] = 12'hfff;
    assign memory[3566] = 12'hfff;
    assign memory[3567] = 12'hfff;
    assign memory[3568] = 12'hfff;
    assign memory[3569] = 12'hfff;
    assign memory[3570] = 12'hfff;
    assign memory[3571] = 12'hfff;
    assign memory[3572] = 12'hfff;
    assign memory[3573] = 12'hfff;
    assign memory[3574] = 12'hfff;
    assign memory[3575] = 12'hfff;
    assign memory[3576] = 12'hfff;
    assign memory[3577] = 12'hfff;
    assign memory[3578] = 12'hfff;
    assign memory[3579] = 12'hfff;
    assign memory[3580] = 12'hfff;
    assign memory[3581] = 12'hfff;
    assign memory[3582] = 12'hfff;
    assign memory[3583] = 12'hfff;
    assign memory[3584] = 12'hfff;
    assign memory[3585] = 12'hfff;
    assign memory[3586] = 12'hfff;
    assign memory[3587] = 12'hfff;
    assign memory[3588] = 12'hfff;
    assign memory[3589] = 12'hfff;
    assign memory[3590] = 12'hfff;
    assign memory[3591] = 12'hfff;
    assign memory[3592] = 12'hfff;
    assign memory[3593] = 12'hfff;
    assign memory[3594] = 12'hfff;
    assign memory[3595] = 12'hfff;
    assign memory[3596] = 12'hfff;
    assign memory[3597] = 12'hfff;
    assign memory[3598] = 12'hfff;
    assign memory[3599] = 12'hfff;
    assign memory[3600] = 12'hfff;
    assign memory[3601] = 12'hfff;
    assign memory[3602] = 12'hfff;
    assign memory[3603] = 12'hfff;
    assign memory[3604] = 12'hfff;
    assign memory[3605] = 12'hfff;
    assign memory[3606] = 12'hfff;
    assign memory[3607] = 12'hfff;
    assign memory[3608] = 12'hfff;
    assign memory[3609] = 12'hfff;
    assign memory[3610] = 12'hfff;
    assign memory[3611] = 12'hfff;
    assign memory[3612] = 12'hfff;
    assign memory[3613] = 12'hfff;
    assign memory[3614] = 12'hfff;
    assign memory[3615] = 12'hfff;
    assign memory[3616] = 12'hfff;
    assign memory[3617] = 12'hfff;
    assign memory[3618] = 12'hfff;
    assign memory[3619] = 12'hfff;
    assign memory[3620] = 12'hfff;
    assign memory[3621] = 12'hfff;
    assign memory[3622] = 12'hfff;
    assign memory[3623] = 12'hfff;
    assign memory[3624] = 12'hfff;
    assign memory[3625] = 12'hfff;
    assign memory[3626] = 12'hfff;
    assign memory[3627] = 12'hfff;
    assign memory[3628] = 12'hfff;
    assign memory[3629] = 12'hfff;
    assign memory[3630] = 12'hfff;
    assign memory[3631] = 12'hfff;
    assign memory[3632] = 12'hfff;
    assign memory[3633] = 12'hfff;
    assign memory[3634] = 12'hfff;
    assign memory[3635] = 12'hfff;
    assign memory[3636] = 12'hfff;
    assign memory[3637] = 12'hfff;
    assign memory[3638] = 12'hfff;
    assign memory[3639] = 12'hfff;
    assign memory[3640] = 12'hfff;
    assign memory[3641] = 12'hfff;
    assign memory[3642] = 12'hfff;
    assign memory[3643] = 12'hfff;
    assign memory[3644] = 12'hfff;
    assign memory[3645] = 12'hfff;
    assign memory[3646] = 12'hfff;
    assign memory[3647] = 12'hfff;
    assign memory[3648] = 12'hfff;
    assign memory[3649] = 12'hfff;
    assign memory[3650] = 12'hfff;
    assign memory[3651] = 12'hfff;
    assign memory[3652] = 12'hfff;
    assign memory[3653] = 12'hfff;
    assign memory[3654] = 12'hfff;
    assign memory[3655] = 12'hfff;
    assign memory[3656] = 12'hfff;
    assign memory[3657] = 12'hfff;
    assign memory[3658] = 12'hfff;
    assign memory[3659] = 12'hfff;
    assign memory[3660] = 12'hfff;
    assign memory[3661] = 12'hfff;
    assign memory[3662] = 12'hfff;
    assign memory[3663] = 12'hfff;
    assign memory[3664] = 12'hfff;
    assign memory[3665] = 12'hfff;
    assign memory[3666] = 12'hfff;
    assign memory[3667] = 12'hfff;
    assign memory[3668] = 12'hfff;
    assign memory[3669] = 12'hfff;
    assign memory[3670] = 12'hfff;
    assign memory[3671] = 12'hfff;
    assign memory[3672] = 12'hfff;
    assign memory[3673] = 12'hfff;
    assign memory[3674] = 12'hfff;
    assign memory[3675] = 12'hfff;
    assign memory[3676] = 12'hfff;
    assign memory[3677] = 12'hfff;
    assign memory[3678] = 12'hfff;
    assign memory[3679] = 12'hfff;
    assign memory[3680] = 12'hfff;
    assign memory[3681] = 12'hfff;
    assign memory[3682] = 12'hfff;
    assign memory[3683] = 12'hfff;
    assign memory[3684] = 12'hfff;
    assign memory[3685] = 12'hfff;
    assign memory[3686] = 12'hfff;
    assign memory[3687] = 12'hfff;
    assign memory[3688] = 12'hfff;
    assign memory[3689] = 12'hfff;
    assign memory[3690] = 12'hfff;
    assign memory[3691] = 12'hfff;
    assign memory[3692] = 12'hfff;
    assign memory[3693] = 12'hfff;
    assign memory[3694] = 12'hfff;
    assign memory[3695] = 12'hfff;
    assign memory[3696] = 12'hfff;
    assign memory[3697] = 12'hfff;
    assign memory[3698] = 12'hfff;
    assign memory[3699] = 12'hfff;
    assign memory[3700] = 12'hfff;
    assign memory[3701] = 12'hfff;
    assign memory[3702] = 12'hfff;
    assign memory[3703] = 12'hfff;
    assign memory[3704] = 12'hfff;
    assign memory[3705] = 12'hfff;
    assign memory[3706] = 12'hfff;
    assign memory[3707] = 12'hfff;
    assign memory[3708] = 12'hfff;
    assign memory[3709] = 12'hfff;
    assign memory[3710] = 12'hfff;
    assign memory[3711] = 12'hfff;
    assign memory[3712] = 12'hfff;
    assign memory[3713] = 12'hfff;
    assign memory[3714] = 12'hfff;
    assign memory[3715] = 12'hfff;
    assign memory[3716] = 12'hfff;
    assign memory[3717] = 12'hfff;
    assign memory[3718] = 12'hfff;
    assign memory[3719] = 12'hfff;
    assign memory[3720] = 12'hfff;
    assign memory[3721] = 12'hfff;
    assign memory[3722] = 12'hfff;
    assign memory[3723] = 12'hfff;
    assign memory[3724] = 12'hfff;
    assign memory[3725] = 12'hfff;
    assign memory[3726] = 12'hfff;
    assign memory[3727] = 12'hfff;
    assign memory[3728] = 12'hfff;
    assign memory[3729] = 12'hfff;
    assign memory[3730] = 12'hfff;
    assign memory[3731] = 12'hfff;
    assign memory[3732] = 12'hfff;
    assign memory[3733] = 12'hfff;
    assign memory[3734] = 12'hfff;
    assign memory[3735] = 12'hfff;
    assign memory[3736] = 12'hfff;
    assign memory[3737] = 12'hfff;
    assign memory[3738] = 12'hfff;
    assign memory[3739] = 12'hfff;
    assign memory[3740] = 12'hfff;
    assign memory[3741] = 12'hfff;
    assign memory[3742] = 12'hfff;
    assign memory[3743] = 12'hfff;
    assign memory[3744] = 12'hfff;
    assign memory[3745] = 12'hfff;
    assign memory[3746] = 12'hfff;
    assign memory[3747] = 12'hfff;
    assign memory[3748] = 12'hfff;
    assign memory[3749] = 12'hfff;
    assign memory[3750] = 12'hfff;
    assign memory[3751] = 12'hfff;
    assign memory[3752] = 12'hfff;
    assign memory[3753] = 12'hfff;
    assign memory[3754] = 12'hfff;
    assign memory[3755] = 12'hfff;
    assign memory[3756] = 12'hfff;
    assign memory[3757] = 12'hfff;
    assign memory[3758] = 12'hfff;
    assign memory[3759] = 12'hfff;
    assign memory[3760] = 12'hfff;
    assign memory[3761] = 12'hfff;
    assign memory[3762] = 12'hfff;
    assign memory[3763] = 12'hfff;
    assign memory[3764] = 12'hfff;
    assign memory[3765] = 12'hfff;
    assign memory[3766] = 12'hfff;
    assign memory[3767] = 12'hfff;
    assign memory[3768] = 12'hfff;
    assign memory[3769] = 12'hfff;
    assign memory[3770] = 12'hfff;
    assign memory[3771] = 12'hfff;
    assign memory[3772] = 12'hfff;
    assign memory[3773] = 12'hfff;
    assign memory[3774] = 12'hfff;
    assign memory[3775] = 12'hfff;
    assign memory[3776] = 12'hfff;
    assign memory[3777] = 12'hfff;
    assign memory[3778] = 12'hfff;
    assign memory[3779] = 12'hfff;
    assign memory[3780] = 12'hfff;
    assign memory[3781] = 12'hfff;
    assign memory[3782] = 12'hfff;
    assign memory[3783] = 12'hfff;
    assign memory[3784] = 12'hfff;
    assign memory[3785] = 12'hfff;
    assign memory[3786] = 12'hfff;
    assign memory[3787] = 12'hfff;
    assign memory[3788] = 12'hfff;
    assign memory[3789] = 12'hfff;
    assign memory[3790] = 12'hfff;
    assign memory[3791] = 12'hfff;
    assign memory[3792] = 12'hfff;
    assign memory[3793] = 12'hfff;
    assign memory[3794] = 12'hfff;
    assign memory[3795] = 12'hfff;
    assign memory[3796] = 12'hfff;
    assign memory[3797] = 12'hfff;
    assign memory[3798] = 12'hfff;
    assign memory[3799] = 12'hfff;
    assign memory[3800] = 12'hfff;
    assign memory[3801] = 12'hfff;
    assign memory[3802] = 12'hfff;
    assign memory[3803] = 12'hfff;
    assign memory[3804] = 12'hfff;
    assign memory[3805] = 12'hfff;
    assign memory[3806] = 12'hfff;
    assign memory[3807] = 12'hfff;
    assign memory[3808] = 12'hfff;
    assign memory[3809] = 12'hfff;
    assign memory[3810] = 12'hfff;
    assign memory[3811] = 12'hfff;
    assign memory[3812] = 12'hfff;
    assign memory[3813] = 12'hfff;
    assign memory[3814] = 12'hfff;
    assign memory[3815] = 12'hfff;
    assign memory[3816] = 12'hfff;
    assign memory[3817] = 12'hfff;
    assign memory[3818] = 12'hfff;
    assign memory[3819] = 12'hfff;
    assign memory[3820] = 12'hfff;
    assign memory[3821] = 12'hfff;
    assign memory[3822] = 12'hfff;
    assign memory[3823] = 12'hfff;
    assign memory[3824] = 12'hfff;
    assign memory[3825] = 12'hfff;
    assign memory[3826] = 12'hfff;
    assign memory[3827] = 12'hfff;
    assign memory[3828] = 12'hfff;
    assign memory[3829] = 12'hfff;
    assign memory[3830] = 12'hfff;
    assign memory[3831] = 12'hfff;
    assign memory[3832] = 12'hfff;
    assign memory[3833] = 12'hfff;
    assign memory[3834] = 12'hfff;
    assign memory[3835] = 12'hfff;
    assign memory[3836] = 12'hfff;
    assign memory[3837] = 12'hfff;
    assign memory[3838] = 12'hfff;
    assign memory[3839] = 12'hfff;
    assign memory[3840] = 12'hfff;
    assign memory[3841] = 12'hfff;
    assign memory[3842] = 12'hfff;
    assign memory[3843] = 12'hfff;
    assign memory[3844] = 12'hfff;
    assign memory[3845] = 12'hfff;
    assign memory[3846] = 12'hfff;
    assign memory[3847] = 12'hfff;
    assign memory[3848] = 12'hfff;
    assign memory[3849] = 12'hfff;
    assign memory[3850] = 12'hfff;
    assign memory[3851] = 12'hfff;
    assign memory[3852] = 12'hfff;
    assign memory[3853] = 12'hfff;
    assign memory[3854] = 12'hfff;
    assign memory[3855] = 12'hfff;
    assign memory[3856] = 12'hfff;
    assign memory[3857] = 12'hfff;
    assign memory[3858] = 12'hfff;
    assign memory[3859] = 12'hfff;
    assign memory[3860] = 12'hfff;
    assign memory[3861] = 12'hfff;
    assign memory[3862] = 12'hfff;
    assign memory[3863] = 12'hfff;
    assign memory[3864] = 12'hfff;
    assign memory[3865] = 12'hfff;
    assign memory[3866] = 12'hfff;
    assign memory[3867] = 12'hfff;
    assign memory[3868] = 12'hfff;
    assign memory[3869] = 12'hfff;
    assign memory[3870] = 12'hfff;
    assign memory[3871] = 12'hfff;
    assign memory[3872] = 12'hfff;
    assign memory[3873] = 12'hfff;
    assign memory[3874] = 12'hfff;
    assign memory[3875] = 12'hfff;
    assign memory[3876] = 12'hfff;
    assign memory[3877] = 12'hfff;
    assign memory[3878] = 12'hfff;
    assign memory[3879] = 12'hfff;
    assign memory[3880] = 12'hfff;
    assign memory[3881] = 12'hfff;
    assign memory[3882] = 12'hfff;
    assign memory[3883] = 12'hfff;
    assign memory[3884] = 12'hfff;
    assign memory[3885] = 12'hfff;
    assign memory[3886] = 12'hfff;
    assign memory[3887] = 12'hfff;
    assign memory[3888] = 12'hfff;
    assign memory[3889] = 12'hfff;
    assign memory[3890] = 12'hfff;
    assign memory[3891] = 12'hfff;
    assign memory[3892] = 12'hfff;
    assign memory[3893] = 12'hfff;
    assign memory[3894] = 12'hfff;
    assign memory[3895] = 12'hfff;
    assign memory[3896] = 12'hfff;
    assign memory[3897] = 12'hfff;
    assign memory[3898] = 12'hfff;
    assign memory[3899] = 12'hfff;
    assign memory[3900] = 12'hfff;
    assign memory[3901] = 12'hfff;
    assign memory[3902] = 12'hfff;
    assign memory[3903] = 12'hfff;
    assign memory[3904] = 12'hfff;
    assign memory[3905] = 12'hfff;
    assign memory[3906] = 12'hfff;
    assign memory[3907] = 12'hfff;
    assign memory[3908] = 12'hfff;
    assign memory[3909] = 12'hfff;
    assign memory[3910] = 12'hfff;
    assign memory[3911] = 12'hfff;
    assign memory[3912] = 12'hfff;
    assign memory[3913] = 12'hfff;
    assign memory[3914] = 12'hfff;
    assign memory[3915] = 12'hfff;
    assign memory[3916] = 12'hfff;
    assign memory[3917] = 12'hfff;
    assign memory[3918] = 12'hfff;
    assign memory[3919] = 12'hfff;
    assign memory[3920] = 12'hfff;
    assign memory[3921] = 12'hfff;
    assign memory[3922] = 12'hfff;
    assign memory[3923] = 12'hfff;
    assign memory[3924] = 12'hfff;
    assign memory[3925] = 12'hfff;
    assign memory[3926] = 12'hfff;
    assign memory[3927] = 12'hfff;
    assign memory[3928] = 12'hfff;
    assign memory[3929] = 12'hfff;
    assign memory[3930] = 12'hfff;
    assign memory[3931] = 12'hfff;
    assign memory[3932] = 12'hfff;
    assign memory[3933] = 12'hfff;
    assign memory[3934] = 12'hfff;
    assign memory[3935] = 12'hfff;
    assign memory[3936] = 12'hfff;
    assign memory[3937] = 12'hfff;
    assign memory[3938] = 12'hfff;
    assign memory[3939] = 12'hfff;
    assign memory[3940] = 12'hfff;
    assign memory[3941] = 12'hfff;
    assign memory[3942] = 12'hfff;
    assign memory[3943] = 12'hfff;
    assign memory[3944] = 12'hfff;
    assign memory[3945] = 12'hfff;
    assign memory[3946] = 12'hfff;
    assign memory[3947] = 12'hfff;
    assign memory[3948] = 12'hfff;
    assign memory[3949] = 12'hfff;
    assign memory[3950] = 12'hfff;
    assign memory[3951] = 12'hfff;
    assign memory[3952] = 12'hfff;
    assign memory[3953] = 12'hfff;
    assign memory[3954] = 12'hfff;
    assign memory[3955] = 12'hfff;
    assign memory[3956] = 12'hfff;
    assign memory[3957] = 12'hfff;
    assign memory[3958] = 12'hfff;
    assign memory[3959] = 12'hfff;
    assign memory[3960] = 12'hfff;
    assign memory[3961] = 12'hfff;
    assign memory[3962] = 12'hfff;
    assign memory[3963] = 12'hfff;
    assign memory[3964] = 12'hfff;
    assign memory[3965] = 12'hfff;
    assign memory[3966] = 12'hfff;
    assign memory[3967] = 12'hfff;
    assign memory[3968] = 12'hfff;
    assign memory[3969] = 12'hfff;
    assign memory[3970] = 12'hfff;
    assign memory[3971] = 12'hfff;
    assign memory[3972] = 12'hfff;
    assign memory[3973] = 12'hfff;
    assign memory[3974] = 12'hfff;
    assign memory[3975] = 12'hfff;
    assign memory[3976] = 12'hfff;
    assign memory[3977] = 12'hfff;
    assign memory[3978] = 12'hfff;
    assign memory[3979] = 12'hfff;
    assign memory[3980] = 12'hfff;
    assign memory[3981] = 12'hfff;
    assign memory[3982] = 12'hfff;
    assign memory[3983] = 12'hfff;
    assign memory[3984] = 12'hfff;
    assign memory[3985] = 12'hfff;
    assign memory[3986] = 12'hfff;
    assign memory[3987] = 12'hfff;
    assign memory[3988] = 12'hfff;
    assign memory[3989] = 12'hfff;
    assign memory[3990] = 12'hfff;
    assign memory[3991] = 12'hfff;
    assign memory[3992] = 12'hfff;
    assign memory[3993] = 12'hfff;
    assign memory[3994] = 12'hfff;
    assign memory[3995] = 12'hfff;
    assign memory[3996] = 12'hfff;
    assign memory[3997] = 12'hfff;
    assign memory[3998] = 12'hfff;
    assign memory[3999] = 12'hfff;
    assign memory[4000] = 12'hfff;
    assign memory[4001] = 12'hfff;
    assign memory[4002] = 12'hfff;
    assign memory[4003] = 12'hfff;
    assign memory[4004] = 12'hfff;
    assign memory[4005] = 12'hfff;
    assign memory[4006] = 12'hfff;
    assign memory[4007] = 12'hfff;
    assign memory[4008] = 12'hfff;
    assign memory[4009] = 12'hfff;
    assign memory[4010] = 12'hfff;
    assign memory[4011] = 12'hfff;
    assign memory[4012] = 12'hfff;
    assign memory[4013] = 12'hfff;
    assign memory[4014] = 12'hfff;
    assign memory[4015] = 12'hfff;
    assign memory[4016] = 12'hfff;
    assign memory[4017] = 12'hfff;
    assign memory[4018] = 12'hfff;
    assign memory[4019] = 12'hfff;
    assign memory[4020] = 12'hfff;
    assign memory[4021] = 12'hfff;
    assign memory[4022] = 12'hfff;
    assign memory[4023] = 12'hfff;
    assign memory[4024] = 12'hfff;
    assign memory[4025] = 12'hfff;
    assign memory[4026] = 12'hfff;
    assign memory[4027] = 12'hfff;
    assign memory[4028] = 12'hfff;
    assign memory[4029] = 12'hfff;
    assign memory[4030] = 12'hfff;
    assign memory[4031] = 12'hfff;
    assign memory[4032] = 12'hfff;
    assign memory[4033] = 12'hfff;
    assign memory[4034] = 12'hfff;
    assign memory[4035] = 12'hfff;
    assign memory[4036] = 12'hfff;
    assign memory[4037] = 12'hfff;
    assign memory[4038] = 12'hfff;
    assign memory[4039] = 12'hfff;
    assign memory[4040] = 12'hfff;
    assign memory[4041] = 12'hfff;
    assign memory[4042] = 12'hfff;
    assign memory[4043] = 12'hfff;
    assign memory[4044] = 12'hfff;
    assign memory[4045] = 12'hfff;
    assign memory[4046] = 12'hfff;
    assign memory[4047] = 12'hfff;
    assign memory[4048] = 12'hfff;
    assign memory[4049] = 12'hfff;
    assign memory[4050] = 12'hfff;
    assign memory[4051] = 12'hfff;
    assign memory[4052] = 12'hfff;
    assign memory[4053] = 12'hfff;
    assign memory[4054] = 12'hfff;
    assign memory[4055] = 12'hfff;
    assign memory[4056] = 12'hfff;
    assign memory[4057] = 12'hfff;
    assign memory[4058] = 12'hfff;
    assign memory[4059] = 12'hfff;
    assign memory[4060] = 12'hfff;
    assign memory[4061] = 12'hfff;
    assign memory[4062] = 12'hfff;
    assign memory[4063] = 12'hfff;
    assign memory[4064] = 12'hfff;
    assign memory[4065] = 12'hfff;
    assign memory[4066] = 12'hfff;
    assign memory[4067] = 12'hfff;
    assign memory[4068] = 12'hfff;
    assign memory[4069] = 12'hfff;
    assign memory[4070] = 12'hfff;
    assign memory[4071] = 12'hfff;
    assign memory[4072] = 12'hfff;
    assign memory[4073] = 12'hfff;
    assign memory[4074] = 12'hfff;
    assign memory[4075] = 12'hfff;
    assign memory[4076] = 12'hfff;
    assign memory[4077] = 12'hfff;
    assign memory[4078] = 12'hfff;
    assign memory[4079] = 12'hfff;
    assign memory[4080] = 12'hfff;
    assign memory[4081] = 12'hfff;
    assign memory[4082] = 12'hfff;
    assign memory[4083] = 12'hfff;
    assign memory[4084] = 12'hfff;
    assign memory[4085] = 12'hfff;
    assign memory[4086] = 12'hfff;
    assign memory[4087] = 12'hfff;
    assign memory[4088] = 12'hfff;
    assign memory[4089] = 12'hfff;
    assign memory[4090] = 12'hfff;
    assign memory[4091] = 12'hfff;
    assign memory[4092] = 12'hfff;
    assign memory[4093] = 12'hfff;
    assign memory[4094] = 12'hfff;
    assign memory[4095] = 12'hfff;
    assign memory[4096] = 12'h890;
    assign memory[4097] = 12'h670;
    assign memory[4098] = 12'hbb0;
    assign memory[4099] = 12'hbb0;
    assign memory[4100] = 12'h670;
    assign memory[4101] = 12'hbb0;
    assign memory[4102] = 12'hbb0;
    assign memory[4103] = 12'hbb0;
    assign memory[4104] = 12'h890;
    assign memory[4105] = 12'hbb0;
    assign memory[4106] = 12'h890;
    assign memory[4107] = 12'hbb0;
    assign memory[4108] = 12'hbb0;
    assign memory[4109] = 12'h670;
    assign memory[4110] = 12'hbb0;
    assign memory[4111] = 12'hbb0;
    assign memory[4112] = 12'hbb0;
    assign memory[4113] = 12'hbb0;
    assign memory[4114] = 12'hbb0;
    assign memory[4115] = 12'h890;
    assign memory[4116] = 12'hbb0;
    assign memory[4117] = 12'h890;
    assign memory[4118] = 12'hbb0;
    assign memory[4119] = 12'hbb0;
    assign memory[4120] = 12'hbb0;
    assign memory[4121] = 12'hbb0;
    assign memory[4122] = 12'h890;
    assign memory[4123] = 12'hbb0;
    assign memory[4124] = 12'hbb0;
    assign memory[4125] = 12'hbb0;
    assign memory[4126] = 12'hbb0;
    assign memory[4127] = 12'hbb0;
    assign memory[4128] = 12'h670;
    assign memory[4129] = 12'hbb0;
    assign memory[4130] = 12'hbb0;
    assign memory[4131] = 12'h670;
    assign memory[4132] = 12'hbb0;
    assign memory[4133] = 12'hbb0;
    assign memory[4134] = 12'hbb0;
    assign memory[4135] = 12'hbb0;
    assign memory[4136] = 12'h890;
    assign memory[4137] = 12'hbb0;
    assign memory[4138] = 12'h890;
    assign memory[4139] = 12'h670;
    assign memory[4140] = 12'hbb0;
    assign memory[4141] = 12'h670;
    assign memory[4142] = 12'hbb0;
    assign memory[4143] = 12'hbb0;
    assign memory[4144] = 12'hbb0;
    assign memory[4145] = 12'hbb0;
    assign memory[4146] = 12'h890;
    assign memory[4147] = 12'h670;
    assign memory[4148] = 12'hbb0;
    assign memory[4149] = 12'hbb0;
    assign memory[4150] = 12'hbb0;
    assign memory[4151] = 12'hbb0;
    assign memory[4152] = 12'hbb0;
    assign memory[4153] = 12'h890;
    assign memory[4154] = 12'h670;
    assign memory[4155] = 12'hbb0;
    assign memory[4156] = 12'hbb0;
    assign memory[4157] = 12'h890;
    assign memory[4158] = 12'hbb0;
    assign memory[4159] = 12'hbb0;
    assign memory[4160] = 12'h890;
    assign memory[4161] = 12'hbb0;
    assign memory[4162] = 12'hbb0;
    assign memory[4163] = 12'h670;
    assign memory[4164] = 12'hbb0;
    assign memory[4165] = 12'hbb0;
    assign memory[4166] = 12'h890;
    assign memory[4167] = 12'hbb0;
    assign memory[4168] = 12'hbb0;
    assign memory[4169] = 12'hbb0;
    assign memory[4170] = 12'hbb0;
    assign memory[4171] = 12'h670;
    assign memory[4172] = 12'hbb0;
    assign memory[4173] = 12'hbb0;
    assign memory[4174] = 12'hbb0;
    assign memory[4175] = 12'hbb0;
    assign memory[4176] = 12'hbb0;
    assign memory[4177] = 12'h890;
    assign memory[4178] = 12'hbb0;
    assign memory[4179] = 12'h670;
    assign memory[4180] = 12'hbb0;
    assign memory[4181] = 12'hbb0;
    assign memory[4182] = 12'hbb0;
    assign memory[4183] = 12'hbb0;
    assign memory[4184] = 12'h890;
    assign memory[4185] = 12'hbb0;
    assign memory[4186] = 12'h670;
    assign memory[4187] = 12'hbb0;
    assign memory[4188] = 12'h890;
    assign memory[4189] = 12'hbb0;
    assign memory[4190] = 12'hbb0;
    assign memory[4191] = 12'h670;
    assign memory[4192] = 12'h890;
    assign memory[4193] = 12'hbb0;
    assign memory[4194] = 12'hbb0;
    assign memory[4195] = 12'h890;
    assign memory[4196] = 12'hbb0;
    assign memory[4197] = 12'hbb0;
    assign memory[4198] = 12'h890;
    assign memory[4199] = 12'h670;
    assign memory[4200] = 12'hbb0;
    assign memory[4201] = 12'hbb0;
    assign memory[4202] = 12'hbb0;
    assign memory[4203] = 12'h670;
    assign memory[4204] = 12'hbb0;
    assign memory[4205] = 12'hbb0;
    assign memory[4206] = 12'hbb0;
    assign memory[4207] = 12'hbb0;
    assign memory[4208] = 12'hbb0;
    assign memory[4209] = 12'h890;
    assign memory[4210] = 12'hbb0;
    assign memory[4211] = 12'h670;
    assign memory[4212] = 12'hbb0;
    assign memory[4213] = 12'h670;
    assign memory[4214] = 12'hbb0;
    assign memory[4215] = 12'hbb0;
    assign memory[4216] = 12'h890;
    assign memory[4217] = 12'hbb0;
    assign memory[4218] = 12'h670;
    assign memory[4219] = 12'hbb0;
    assign memory[4220] = 12'h890;
    assign memory[4221] = 12'hbb0;
    assign memory[4222] = 12'hbb0;
    assign memory[4223] = 12'h670;
    assign memory[4224] = 12'h890;
    assign memory[4225] = 12'hbb0;
    assign memory[4226] = 12'h890;
    assign memory[4227] = 12'h670;
    assign memory[4228] = 12'hbb0;
    assign memory[4229] = 12'hbb0;
    assign memory[4230] = 12'h890;
    assign memory[4231] = 12'h670;
    assign memory[4232] = 12'hbb0;
    assign memory[4233] = 12'hbb0;
    assign memory[4234] = 12'hbb0;
    assign memory[4235] = 12'h670;
    assign memory[4236] = 12'h890;
    assign memory[4237] = 12'hbb0;
    assign memory[4238] = 12'hbb0;
    assign memory[4239] = 12'h670;
    assign memory[4240] = 12'hbb0;
    assign memory[4241] = 12'h890;
    assign memory[4242] = 12'hbb0;
    assign memory[4243] = 12'h670;
    assign memory[4244] = 12'hbb0;
    assign memory[4245] = 12'h670;
    assign memory[4246] = 12'hbb0;
    assign memory[4247] = 12'hbb0;
    assign memory[4248] = 12'h890;
    assign memory[4249] = 12'hbb0;
    assign memory[4250] = 12'h670;
    assign memory[4251] = 12'hbb0;
    assign memory[4252] = 12'h890;
    assign memory[4253] = 12'hbb0;
    assign memory[4254] = 12'hbb0;
    assign memory[4255] = 12'h670;
    assign memory[4256] = 12'h890;
    assign memory[4257] = 12'hbb0;
    assign memory[4258] = 12'h890;
    assign memory[4259] = 12'h670;
    assign memory[4260] = 12'hbb0;
    assign memory[4261] = 12'hbb0;
    assign memory[4262] = 12'h890;
    assign memory[4263] = 12'h670;
    assign memory[4264] = 12'hbb0;
    assign memory[4265] = 12'hbb0;
    assign memory[4266] = 12'hbb0;
    assign memory[4267] = 12'hbb0;
    assign memory[4268] = 12'h890;
    assign memory[4269] = 12'hbb0;
    assign memory[4270] = 12'hbb0;
    assign memory[4271] = 12'h670;
    assign memory[4272] = 12'hbb0;
    assign memory[4273] = 12'h890;
    assign memory[4274] = 12'hbb0;
    assign memory[4275] = 12'hbb0;
    assign memory[4276] = 12'h890;
    assign memory[4277] = 12'h670;
    assign memory[4278] = 12'hbb0;
    assign memory[4279] = 12'hbb0;
    assign memory[4280] = 12'h890;
    assign memory[4281] = 12'hbb0;
    assign memory[4282] = 12'hbb0;
    assign memory[4283] = 12'hbb0;
    assign memory[4284] = 12'h890;
    assign memory[4285] = 12'h670;
    assign memory[4286] = 12'hbb0;
    assign memory[4287] = 12'h670;
    assign memory[4288] = 12'h890;
    assign memory[4289] = 12'hbb0;
    assign memory[4290] = 12'h890;
    assign memory[4291] = 12'h670;
    assign memory[4292] = 12'h890;
    assign memory[4293] = 12'hbb0;
    assign memory[4294] = 12'h890;
    assign memory[4295] = 12'h670;
    assign memory[4296] = 12'h890;
    assign memory[4297] = 12'hbb0;
    assign memory[4298] = 12'hbb0;
    assign memory[4299] = 12'hbb0;
    assign memory[4300] = 12'h890;
    assign memory[4301] = 12'hbb0;
    assign memory[4302] = 12'hbb0;
    assign memory[4303] = 12'h670;
    assign memory[4304] = 12'hbb0;
    assign memory[4305] = 12'h890;
    assign memory[4306] = 12'hbb0;
    assign memory[4307] = 12'hbb0;
    assign memory[4308] = 12'h890;
    assign memory[4309] = 12'h670;
    assign memory[4310] = 12'hbb0;
    assign memory[4311] = 12'h670;
    assign memory[4312] = 12'h890;
    assign memory[4313] = 12'hbb0;
    assign memory[4314] = 12'hbb0;
    assign memory[4315] = 12'hbb0;
    assign memory[4316] = 12'h890;
    assign memory[4317] = 12'h670;
    assign memory[4318] = 12'h890;
    assign memory[4319] = 12'hbb0;
    assign memory[4320] = 12'hbb0;
    assign memory[4321] = 12'hbb0;
    assign memory[4322] = 12'h890;
    assign memory[4323] = 12'hbb0;
    assign memory[4324] = 12'h890;
    assign memory[4325] = 12'hbb0;
    assign memory[4326] = 12'hbb0;
    assign memory[4327] = 12'h670;
    assign memory[4328] = 12'h890;
    assign memory[4329] = 12'hbb0;
    assign memory[4330] = 12'hbb0;
    assign memory[4331] = 12'hbb0;
    assign memory[4332] = 12'h890;
    assign memory[4333] = 12'hbb0;
    assign memory[4334] = 12'h890;
    assign memory[4335] = 12'h670;
    assign memory[4336] = 12'hbb0;
    assign memory[4337] = 12'hbb0;
    assign memory[4338] = 12'hbb0;
    assign memory[4339] = 12'hbb0;
    assign memory[4340] = 12'h890;
    assign memory[4341] = 12'h670;
    assign memory[4342] = 12'hbb0;
    assign memory[4343] = 12'h670;
    assign memory[4344] = 12'hbb0;
    assign memory[4345] = 12'hbb0;
    assign memory[4346] = 12'hbb0;
    assign memory[4347] = 12'h670;
    assign memory[4348] = 12'hbb0;
    assign memory[4349] = 12'h670;
    assign memory[4350] = 12'h890;
    assign memory[4351] = 12'hbb0;
    assign memory[4352] = 12'hbb0;
    assign memory[4353] = 12'hbb0;
    assign memory[4354] = 12'h890;
    assign memory[4355] = 12'hbb0;
    assign memory[4356] = 12'h890;
    assign memory[4357] = 12'hbb0;
    assign memory[4358] = 12'hbb0;
    assign memory[4359] = 12'h670;
    assign memory[4360] = 12'h890;
    assign memory[4361] = 12'h670;
    assign memory[4362] = 12'hbb0;
    assign memory[4363] = 12'hbb0;
    assign memory[4364] = 12'h890;
    assign memory[4365] = 12'hbb0;
    assign memory[4366] = 12'h890;
    assign memory[4367] = 12'h670;
    assign memory[4368] = 12'hbb0;
    assign memory[4369] = 12'hbb0;
    assign memory[4370] = 12'hbb0;
    assign memory[4371] = 12'h670;
    assign memory[4372] = 12'h890;
    assign memory[4373] = 12'hbb0;
    assign memory[4374] = 12'hbb0;
    assign memory[4375] = 12'h670;
    assign memory[4376] = 12'hbb0;
    assign memory[4377] = 12'hbb0;
    assign memory[4378] = 12'hbb0;
    assign memory[4379] = 12'h670;
    assign memory[4380] = 12'hbb0;
    assign memory[4381] = 12'h670;
    assign memory[4382] = 12'h890;
    assign memory[4383] = 12'h670;
    assign memory[4384] = 12'hbb0;
    assign memory[4385] = 12'h670;
    assign memory[4386] = 12'hbb0;
    assign memory[4387] = 12'hbb0;
    assign memory[4388] = 12'h890;
    assign memory[4389] = 12'hbb0;
    assign memory[4390] = 12'hbb0;
    assign memory[4391] = 12'hbb0;
    assign memory[4392] = 12'h890;
    assign memory[4393] = 12'h670;
    assign memory[4394] = 12'hbb0;
    assign memory[4395] = 12'hbb0;
    assign memory[4396] = 12'h890;
    assign memory[4397] = 12'hbb0;
    assign memory[4398] = 12'h890;
    assign memory[4399] = 12'h670;
    assign memory[4400] = 12'hbb0;
    assign memory[4401] = 12'hbb0;
    assign memory[4402] = 12'hbb0;
    assign memory[4403] = 12'h670;
    assign memory[4404] = 12'h890;
    assign memory[4405] = 12'hbb0;
    assign memory[4406] = 12'hbb0;
    assign memory[4407] = 12'h670;
    assign memory[4408] = 12'hbb0;
    assign memory[4409] = 12'h780;
    assign memory[4410] = 12'h890;
    assign memory[4411] = 12'h670;
    assign memory[4412] = 12'hbb0;
    assign memory[4413] = 12'hbb0;
    assign memory[4414] = 12'h890;
    assign memory[4415] = 12'h670;
    assign memory[4416] = 12'hbb0;
    assign memory[4417] = 12'h670;
    assign memory[4418] = 12'hbb0;
    assign memory[4419] = 12'hbb0;
    assign memory[4420] = 12'h890;
    assign memory[4421] = 12'hbb0;
    assign memory[4422] = 12'h890;
    assign memory[4423] = 12'hbb0;
    assign memory[4424] = 12'hbb0;
    assign memory[4425] = 12'h670;
    assign memory[4426] = 12'hbb0;
    assign memory[4427] = 12'h890;
    assign memory[4428] = 12'hbb0;
    assign memory[4429] = 12'hbb0;
    assign memory[4430] = 12'h890;
    assign memory[4431] = 12'hbb0;
    assign memory[4432] = 12'hbb0;
    assign memory[4433] = 12'hbb0;
    assign memory[4434] = 12'h890;
    assign memory[4435] = 12'h670;
    assign memory[4436] = 12'hbb0;
    assign memory[4437] = 12'hbb0;
    assign memory[4438] = 12'hbb0;
    assign memory[4439] = 12'h670;
    assign memory[4440] = 12'h780;
    assign memory[4441] = 12'h670;
    assign memory[4442] = 12'h890;
    assign memory[4443] = 12'h670;
    assign memory[4444] = 12'hbb0;
    assign memory[4445] = 12'hbb0;
    assign memory[4446] = 12'h890;
    assign memory[4447] = 12'h670;
    assign memory[4448] = 12'hbb0;
    assign memory[4449] = 12'h670;
    assign memory[4450] = 12'hbb0;
    assign memory[4451] = 12'hbb0;
    assign memory[4452] = 12'h890;
    assign memory[4453] = 12'hbb0;
    assign memory[4454] = 12'h890;
    assign memory[4455] = 12'hbb0;
    assign memory[4456] = 12'hbb0;
    assign memory[4457] = 12'h670;
    assign memory[4458] = 12'hbb0;
    assign memory[4459] = 12'h890;
    assign memory[4460] = 12'hbb0;
    assign memory[4461] = 12'hbb0;
    assign memory[4462] = 12'h890;
    assign memory[4463] = 12'hbb0;
    assign memory[4464] = 12'hbb0;
    assign memory[4465] = 12'hbb0;
    assign memory[4466] = 12'h780;
    assign memory[4467] = 12'h670;
    assign memory[4468] = 12'hbb0;
    assign memory[4469] = 12'hbb0;
    assign memory[4470] = 12'hbb0;
    assign memory[4471] = 12'h780;
    assign memory[4472] = 12'hbb0;
    assign memory[4473] = 12'h670;
    assign memory[4474] = 12'h890;
    assign memory[4475] = 12'h670;
    assign memory[4476] = 12'hbb0;
    assign memory[4477] = 12'h670;
    assign memory[4478] = 12'h890;
    assign memory[4479] = 12'h670;
    assign memory[4480] = 12'hbb0;
    assign memory[4481] = 12'h670;
    assign memory[4482] = 12'hbb0;
    assign memory[4483] = 12'hbb0;
    assign memory[4484] = 12'h890;
    assign memory[4485] = 12'hbb0;
    assign memory[4486] = 12'h890;
    assign memory[4487] = 12'hbb0;
    assign memory[4488] = 12'hbb0;
    assign memory[4489] = 12'h670;
    assign memory[4490] = 12'hbb0;
    assign memory[4491] = 12'h890;
    assign memory[4492] = 12'hbb0;
    assign memory[4493] = 12'hbb0;
    assign memory[4494] = 12'h890;
    assign memory[4495] = 12'hbb0;
    assign memory[4496] = 12'hbb0;
    assign memory[4497] = 12'h780;
    assign memory[4498] = 12'h890;
    assign memory[4499] = 12'h670;
    assign memory[4500] = 12'hbb0;
    assign memory[4501] = 12'hbb0;
    assign memory[4502] = 12'hbb0;
    assign memory[4503] = 12'h780;
    assign memory[4504] = 12'hbb0;
    assign memory[4505] = 12'h670;
    assign memory[4506] = 12'h890;
    assign memory[4507] = 12'h670;
    assign memory[4508] = 12'hbb0;
    assign memory[4509] = 12'h670;
    assign memory[4510] = 12'hbb0;
    assign memory[4511] = 12'h670;
    assign memory[4512] = 12'h890;
    assign memory[4513] = 12'h670;
    assign memory[4514] = 12'hbb0;
    assign memory[4515] = 12'hbb0;
    assign memory[4516] = 12'hbb0;
    assign memory[4517] = 12'hbb0;
    assign memory[4518] = 12'h890;
    assign memory[4519] = 12'hbb0;
    assign memory[4520] = 12'hbb0;
    assign memory[4521] = 12'hbb0;
    assign memory[4522] = 12'hbb0;
    assign memory[4523] = 12'h890;
    assign memory[4524] = 12'h670;
    assign memory[4525] = 12'hbb0;
    assign memory[4526] = 12'h890;
    assign memory[4527] = 12'hbb0;
    assign memory[4528] = 12'h780;
    assign memory[4529] = 12'hbb0;
    assign memory[4530] = 12'h890;
    assign memory[4531] = 12'hbb0;
    assign memory[4532] = 12'hbb0;
    assign memory[4533] = 12'h670;
    assign memory[4534] = 12'hbb0;
    assign memory[4535] = 12'h780;
    assign memory[4536] = 12'hbb0;
    assign memory[4537] = 12'h670;
    assign memory[4538] = 12'h890;
    assign memory[4539] = 12'hbb0;
    assign memory[4540] = 12'hbb0;
    assign memory[4541] = 12'h670;
    assign memory[4542] = 12'hbb0;
    assign memory[4543] = 12'hbb0;
    assign memory[4544] = 12'h890;
    assign memory[4545] = 12'h670;
    assign memory[4546] = 12'hbb0;
    assign memory[4547] = 12'hbb0;
    assign memory[4548] = 12'hbb0;
    assign memory[4549] = 12'h670;
    assign memory[4550] = 12'h890;
    assign memory[4551] = 12'hbb0;
    assign memory[4552] = 12'hbb0;
    assign memory[4553] = 12'hbb0;
    assign memory[4554] = 12'hbb0;
    assign memory[4555] = 12'h890;
    assign memory[4556] = 12'h670;
    assign memory[4557] = 12'hbb0;
    assign memory[4558] = 12'hbb0;
    assign memory[4559] = 12'hbb0;
    assign memory[4560] = 12'h780;
    assign memory[4561] = 12'hbb0;
    assign memory[4562] = 12'h890;
    assign memory[4563] = 12'hbb0;
    assign memory[4564] = 12'hbb0;
    assign memory[4565] = 12'h670;
    assign memory[4566] = 12'hbb0;
    assign memory[4567] = 12'h780;
    assign memory[4568] = 12'hbb0;
    assign memory[4569] = 12'h670;
    assign memory[4570] = 12'hbb0;
    assign memory[4571] = 12'hbb0;
    assign memory[4572] = 12'hbb0;
    assign memory[4573] = 12'h670;
    assign memory[4574] = 12'hbb0;
    assign memory[4575] = 12'hbb0;
    assign memory[4576] = 12'h890;
    assign memory[4577] = 12'hbb0;
    assign memory[4578] = 12'hbb0;
    assign memory[4579] = 12'hbb0;
    assign memory[4580] = 12'hbb0;
    assign memory[4581] = 12'h670;
    assign memory[4582] = 12'hbb0;
    assign memory[4583] = 12'hbb0;
    assign memory[4584] = 12'h890;
    assign memory[4585] = 12'hbb0;
    assign memory[4586] = 12'hbb0;
    assign memory[4587] = 12'hbb0;
    assign memory[4588] = 12'h670;
    assign memory[4589] = 12'hbb0;
    assign memory[4590] = 12'hbb0;
    assign memory[4591] = 12'hbb0;
    assign memory[4592] = 12'h780;
    assign memory[4593] = 12'hbb0;
    assign memory[4594] = 12'hbb0;
    assign memory[4595] = 12'hbb0;
    assign memory[4596] = 12'h890;
    assign memory[4597] = 12'h670;
    assign memory[4598] = 12'hbb0;
    assign memory[4599] = 12'h780;
    assign memory[4600] = 12'hbb0;
    assign memory[4601] = 12'hbb0;
    assign memory[4602] = 12'hbb0;
    assign memory[4603] = 12'hbb0;
    assign memory[4604] = 12'hbb0;
    assign memory[4605] = 12'h670;
    assign memory[4606] = 12'hbb0;
    assign memory[4607] = 12'hbb0;
    assign memory[4608] = 12'h890;
    assign memory[4609] = 12'hbb0;
    assign memory[4610] = 12'hbb0;
    assign memory[4611] = 12'h890;
    assign memory[4612] = 12'hbb0;
    assign memory[4613] = 12'h670;
    assign memory[4614] = 12'hbb0;
    assign memory[4615] = 12'h890;
    assign memory[4616] = 12'hbb0;
    assign memory[4617] = 12'hbb0;
    assign memory[4618] = 12'hbb0;
    assign memory[4619] = 12'hbb0;
    assign memory[4620] = 12'h670;
    assign memory[4621] = 12'hbb0;
    assign memory[4622] = 12'hbb0;
    assign memory[4623] = 12'hbb0;
    assign memory[4624] = 12'h780;
    assign memory[4625] = 12'h670;
    assign memory[4626] = 12'hbb0;
    assign memory[4627] = 12'hbb0;
    assign memory[4628] = 12'h890;
    assign memory[4629] = 12'h670;
    assign memory[4630] = 12'hbb0;
    assign memory[4631] = 12'hbb0;
    assign memory[4632] = 12'h890;
    assign memory[4633] = 12'hbb0;
    assign memory[4634] = 12'hbb0;
    assign memory[4635] = 12'hbb0;
    assign memory[4636] = 12'h890;
    assign memory[4637] = 12'h670;
    assign memory[4638] = 12'hbb0;
    assign memory[4639] = 12'hbb0;
    assign memory[4640] = 12'h890;
    assign memory[4641] = 12'hbb0;
    assign memory[4642] = 12'h670;
    assign memory[4643] = 12'h890;
    assign memory[4644] = 12'hbb0;
    assign memory[4645] = 12'h670;
    assign memory[4646] = 12'hbb0;
    assign memory[4647] = 12'h890;
    assign memory[4648] = 12'hbb0;
    assign memory[4649] = 12'h890;
    assign memory[4650] = 12'hbb0;
    assign memory[4651] = 12'hbb0;
    assign memory[4652] = 12'h670;
    assign memory[4653] = 12'hbb0;
    assign memory[4654] = 12'hbb0;
    assign memory[4655] = 12'hbb0;
    assign memory[4656] = 12'h780;
    assign memory[4657] = 12'h670;
    assign memory[4658] = 12'hbb0;
    assign memory[4659] = 12'hbb0;
    assign memory[4660] = 12'h890;
    assign memory[4661] = 12'h670;
    assign memory[4662] = 12'hbb0;
    assign memory[4663] = 12'hbb0;
    assign memory[4664] = 12'h890;
    assign memory[4665] = 12'hbb0;
    assign memory[4666] = 12'h670;
    assign memory[4667] = 12'hbb0;
    assign memory[4668] = 12'h890;
    assign memory[4669] = 12'hbb0;
    assign memory[4670] = 12'hbb0;
    assign memory[4671] = 12'hbb0;
    assign memory[4672] = 12'h890;
    assign memory[4673] = 12'hbb0;
    assign memory[4674] = 12'h670;
    assign memory[4675] = 12'h890;
    assign memory[4676] = 12'hbb0;
    assign memory[4677] = 12'h670;
    assign memory[4678] = 12'hbb0;
    assign memory[4679] = 12'h890;
    assign memory[4680] = 12'hbb0;
    assign memory[4681] = 12'h890;
    assign memory[4682] = 12'hbb0;
    assign memory[4683] = 12'hbb0;
    assign memory[4684] = 12'hbb0;
    assign memory[4685] = 12'hbb0;
    assign memory[4686] = 12'h780;
    assign memory[4687] = 12'hbb0;
    assign memory[4688] = 12'h780;
    assign memory[4689] = 12'h670;
    assign memory[4690] = 12'hbb0;
    assign memory[4691] = 12'hbb0;
    assign memory[4692] = 12'h890;
    assign memory[4693] = 12'hbb0;
    assign memory[4694] = 12'hbb0;
    assign memory[4695] = 12'hbb0;
    assign memory[4696] = 12'h890;
    assign memory[4697] = 12'hbb0;
    assign memory[4698] = 12'h670;
    assign memory[4699] = 12'hbb0;
    assign memory[4700] = 12'h890;
    assign memory[4701] = 12'hbb0;
    assign memory[4702] = 12'hbb0;
    assign memory[4703] = 12'hbb0;
    assign memory[4704] = 12'hbb0;
    assign memory[4705] = 12'hbb0;
    assign memory[4706] = 12'h670;
    assign memory[4707] = 12'h890;
    assign memory[4708] = 12'hbb0;
    assign memory[4709] = 12'h670;
    assign memory[4710] = 12'hbb0;
    assign memory[4711] = 12'h890;
    assign memory[4712] = 12'hbb0;
    assign memory[4713] = 12'h890;
    assign memory[4714] = 12'hbb0;
    assign memory[4715] = 12'hbb0;
    assign memory[4716] = 12'hbb0;
    assign memory[4717] = 12'h780;
    assign memory[4718] = 12'hbb0;
    assign memory[4719] = 12'h890;
    assign memory[4720] = 12'hbb0;
    assign memory[4721] = 12'h670;
    assign memory[4722] = 12'hbb0;
    assign memory[4723] = 12'hbb0;
    assign memory[4724] = 12'h890;
    assign memory[4725] = 12'hbb0;
    assign memory[4726] = 12'hbb0;
    assign memory[4727] = 12'hbb0;
    assign memory[4728] = 12'h890;
    assign memory[4729] = 12'hbb0;
    assign memory[4730] = 12'h670;
    assign memory[4731] = 12'hbb0;
    assign memory[4732] = 12'h890;
    assign memory[4733] = 12'h670;
    assign memory[4734] = 12'hbb0;
    assign memory[4735] = 12'hbb0;
    assign memory[4736] = 12'hbb0;
    assign memory[4737] = 12'hbb0;
    assign memory[4738] = 12'h670;
    assign memory[4739] = 12'h890;
    assign memory[4740] = 12'hbb0;
    assign memory[4741] = 12'hbb0;
    assign memory[4742] = 12'hbb0;
    assign memory[4743] = 12'h890;
    assign memory[4744] = 12'hbb0;
    assign memory[4745] = 12'h890;
    assign memory[4746] = 12'h670;
    assign memory[4747] = 12'h890;
    assign memory[4748] = 12'h780;
    assign memory[4749] = 12'hbb0;
    assign memory[4750] = 12'hbb0;
    assign memory[4751] = 12'h890;
    assign memory[4752] = 12'hbb0;
    assign memory[4753] = 12'h670;
    assign memory[4754] = 12'hbb0;
    assign memory[4755] = 12'hbb0;
    assign memory[4756] = 12'hbb0;
    assign memory[4757] = 12'hbb0;
    assign memory[4758] = 12'hbb0;
    assign memory[4759] = 12'h670;
    assign memory[4760] = 12'h890;
    assign memory[4761] = 12'hbb0;
    assign memory[4762] = 12'h670;
    assign memory[4763] = 12'hbb0;
    assign memory[4764] = 12'h890;
    assign memory[4765] = 12'h670;
    assign memory[4766] = 12'hbb0;
    assign memory[4767] = 12'hbb0;
    assign memory[4768] = 12'hbb0;
    assign memory[4769] = 12'h890;
    assign memory[4770] = 12'h670;
    assign memory[4771] = 12'h890;
    assign memory[4772] = 12'hbb0;
    assign memory[4773] = 12'hbb0;
    assign memory[4774] = 12'hbb0;
    assign memory[4775] = 12'h890;
    assign memory[4776] = 12'hbb0;
    assign memory[4777] = 12'h890;
    assign memory[4778] = 12'h670;
    assign memory[4779] = 12'h890;
    assign memory[4780] = 12'h780;
    assign memory[4781] = 12'hbb0;
    assign memory[4782] = 12'h670;
    assign memory[4783] = 12'h890;
    assign memory[4784] = 12'hbb0;
    assign memory[4785] = 12'h670;
    assign memory[4786] = 12'hbb0;
    assign memory[4787] = 12'hbb0;
    assign memory[4788] = 12'h670;
    assign memory[4789] = 12'hbb0;
    assign memory[4790] = 12'h890;
    assign memory[4791] = 12'h670;
    assign memory[4792] = 12'hbb0;
    assign memory[4793] = 12'hbb0;
    assign memory[4794] = 12'h670;
    assign memory[4795] = 12'hbb0;
    assign memory[4796] = 12'hbb0;
    assign memory[4797] = 12'h670;
    assign memory[4798] = 12'hbb0;
    assign memory[4799] = 12'h670;
    assign memory[4800] = 12'hbb0;
    assign memory[4801] = 12'h890;
    assign memory[4802] = 12'hbb0;
    assign memory[4803] = 12'hbb0;
    assign memory[4804] = 12'hbb0;
    assign memory[4805] = 12'hbb0;
    assign memory[4806] = 12'hbb0;
    assign memory[4807] = 12'hbb0;
    assign memory[4808] = 12'hbb0;
    assign memory[4809] = 12'hbb0;
    assign memory[4810] = 12'h670;
    assign memory[4811] = 12'h890;
    assign memory[4812] = 12'h780;
    assign memory[4813] = 12'hbb0;
    assign memory[4814] = 12'h670;
    assign memory[4815] = 12'h890;
    assign memory[4816] = 12'hbb0;
    assign memory[4817] = 12'h670;
    assign memory[4818] = 12'h890;
    assign memory[4819] = 12'hbb0;
    assign memory[4820] = 12'h670;
    assign memory[4821] = 12'hbb0;
    assign memory[4822] = 12'h890;
    assign memory[4823] = 12'h670;
    assign memory[4824] = 12'hbb0;
    assign memory[4825] = 12'hbb0;
    assign memory[4826] = 12'hbb0;
    assign memory[4827] = 12'hbb0;
    assign memory[4828] = 12'hbb0;
    assign memory[4829] = 12'h670;
    assign memory[4830] = 12'hbb0;
    assign memory[4831] = 12'h670;
    assign memory[4832] = 12'hbb0;
    assign memory[4833] = 12'h890;
    assign memory[4834] = 12'hbb0;
    assign memory[4835] = 12'hbb0;
    assign memory[4836] = 12'hbb0;
    assign memory[4837] = 12'hbb0;
    assign memory[4838] = 12'h890;
    assign memory[4839] = 12'hbb0;
    assign memory[4840] = 12'hbb0;
    assign memory[4841] = 12'hbb0;
    assign memory[4842] = 12'h670;
    assign memory[4843] = 12'h890;
    assign memory[4844] = 12'h780;
    assign memory[4845] = 12'hbb0;
    assign memory[4846] = 12'h670;
    assign memory[4847] = 12'h890;
    assign memory[4848] = 12'hbb0;
    assign memory[4849] = 12'hbb0;
    assign memory[4850] = 12'h890;
    assign memory[4851] = 12'hbb0;
    assign memory[4852] = 12'h670;
    assign memory[4853] = 12'hbb0;
    assign memory[4854] = 12'h890;
    assign memory[4855] = 12'h670;
    assign memory[4856] = 12'hbb0;
    assign memory[4857] = 12'hbb0;
    assign memory[4858] = 12'hbb0;
    assign memory[4859] = 12'hbb0;
    assign memory[4860] = 12'hbb0;
    assign memory[4861] = 12'h670;
    assign memory[4862] = 12'hbb0;
    assign memory[4863] = 12'h670;
    assign memory[4864] = 12'hbb0;
    assign memory[4865] = 12'h890;
    assign memory[4866] = 12'hbb0;
    assign memory[4867] = 12'hbb0;
    assign memory[4868] = 12'hbb0;
    assign memory[4869] = 12'h890;
    assign memory[4870] = 12'hbb0;
    assign memory[4871] = 12'h670;
    assign memory[4872] = 12'hbb0;
    assign memory[4873] = 12'hbb0;
    assign memory[4874] = 12'h670;
    assign memory[4875] = 12'h890;
    assign memory[4876] = 12'h780;
    assign memory[4877] = 12'hbb0;
    assign memory[4878] = 12'h670;
    assign memory[4879] = 12'h890;
    assign memory[4880] = 12'hbb0;
    assign memory[4881] = 12'hbb0;
    assign memory[4882] = 12'h890;
    assign memory[4883] = 12'hbb0;
    assign memory[4884] = 12'h670;
    assign memory[4885] = 12'hbb0;
    assign memory[4886] = 12'h890;
    assign memory[4887] = 12'h670;
    assign memory[4888] = 12'hbb0;
    assign memory[4889] = 12'hbb0;
    assign memory[4890] = 12'h780;
    assign memory[4891] = 12'h670;
    assign memory[4892] = 12'hbb0;
    assign memory[4893] = 12'hbb0;
    assign memory[4894] = 12'hbb0;
    assign memory[4895] = 12'h670;
    assign memory[4896] = 12'hbb0;
    assign memory[4897] = 12'h890;
    assign memory[4898] = 12'hbb0;
    assign memory[4899] = 12'hbb0;
    assign memory[4900] = 12'hbb0;
    assign memory[4901] = 12'h890;
    assign memory[4902] = 12'hbb0;
    assign memory[4903] = 12'h670;
    assign memory[4904] = 12'hbb0;
    assign memory[4905] = 12'h890;
    assign memory[4906] = 12'h670;
    assign memory[4907] = 12'hbb0;
    assign memory[4908] = 12'h780;
    assign memory[4909] = 12'hbb0;
    assign memory[4910] = 12'h670;
    assign memory[4911] = 12'hbb0;
    assign memory[4912] = 12'hbb0;
    assign memory[4913] = 12'hbb0;
    assign memory[4914] = 12'h890;
    assign memory[4915] = 12'hbb0;
    assign memory[4916] = 12'h670;
    assign memory[4917] = 12'hbb0;
    assign memory[4918] = 12'h890;
    assign memory[4919] = 12'h670;
    assign memory[4920] = 12'hbb0;
    assign memory[4921] = 12'h780;
    assign memory[4922] = 12'h890;
    assign memory[4923] = 12'h670;
    assign memory[4924] = 12'hbb0;
    assign memory[4925] = 12'hbb0;
    assign memory[4926] = 12'hbb0;
    assign memory[4927] = 12'h670;
    assign memory[4928] = 12'hbb0;
    assign memory[4929] = 12'hbb0;
    assign memory[4930] = 12'hbb0;
    assign memory[4931] = 12'h890;
    assign memory[4932] = 12'hbb0;
    assign memory[4933] = 12'h890;
    assign memory[4934] = 12'hbb0;
    assign memory[4935] = 12'h670;
    assign memory[4936] = 12'h890;
    assign memory[4937] = 12'hbb0;
    assign memory[4938] = 12'hbb0;
    assign memory[4939] = 12'hbb0;
    assign memory[4940] = 12'hbb0;
    assign memory[4941] = 12'h890;
    assign memory[4942] = 12'hbb0;
    assign memory[4943] = 12'hbb0;
    assign memory[4944] = 12'hbb0;
    assign memory[4945] = 12'hbb0;
    assign memory[4946] = 12'hbb0;
    assign memory[4947] = 12'hbb0;
    assign memory[4948] = 12'h670;
    assign memory[4949] = 12'hbb0;
    assign memory[4950] = 12'hbb0;
    assign memory[4951] = 12'hbb0;
    assign memory[4952] = 12'h780;
    assign memory[4953] = 12'hbb0;
    assign memory[4954] = 12'h890;
    assign memory[4955] = 12'h670;
    assign memory[4956] = 12'hbb0;
    assign memory[4957] = 12'hbb0;
    assign memory[4958] = 12'hbb0;
    assign memory[4959] = 12'h670;
    assign memory[4960] = 12'hbb0;
    assign memory[4961] = 12'hbb0;
    assign memory[4962] = 12'h890;
    assign memory[4963] = 12'hbb0;
    assign memory[4964] = 12'hbb0;
    assign memory[4965] = 12'h890;
    assign memory[4966] = 12'hbb0;
    assign memory[4967] = 12'h670;
    assign memory[4968] = 12'h890;
    assign memory[4969] = 12'hbb0;
    assign memory[4970] = 12'hbb0;
    assign memory[4971] = 12'hbb0;
    assign memory[4972] = 12'h890;
    assign memory[4973] = 12'hbb0;
    assign memory[4974] = 12'hbb0;
    assign memory[4975] = 12'hbb0;
    assign memory[4976] = 12'hbb0;
    assign memory[4977] = 12'hbb0;
    assign memory[4978] = 12'hbb0;
    assign memory[4979] = 12'hbb0;
    assign memory[4980] = 12'hbb0;
    assign memory[4981] = 12'hbb0;
    assign memory[4982] = 12'hbb0;
    assign memory[4983] = 12'h890;
    assign memory[4984] = 12'h780;
    assign memory[4985] = 12'hbb0;
    assign memory[4986] = 12'h890;
    assign memory[4987] = 12'h670;
    assign memory[4988] = 12'hbb0;
    assign memory[4989] = 12'hbb0;
    assign memory[4990] = 12'hbb0;
    assign memory[4991] = 12'hbb0;
    assign memory[4992] = 12'hbb0;
    assign memory[4993] = 12'hbb0;
    assign memory[4994] = 12'h890;
    assign memory[4995] = 12'hbb0;
    assign memory[4996] = 12'h670;
    assign memory[4997] = 12'h890;
    assign memory[4998] = 12'hbb0;
    assign memory[4999] = 12'h670;
    assign memory[5000] = 12'h890;
    assign memory[5001] = 12'hbb0;
    assign memory[5002] = 12'hbb0;
    assign memory[5003] = 12'hbb0;
    assign memory[5004] = 12'h890;
    assign memory[5005] = 12'hbb0;
    assign memory[5006] = 12'hbb0;
    assign memory[5007] = 12'h670;
    assign memory[5008] = 12'hbb0;
    assign memory[5009] = 12'hbb0;
    assign memory[5010] = 12'h670;
    assign memory[5011] = 12'hbb0;
    assign memory[5012] = 12'hbb0;
    assign memory[5013] = 12'hbb0;
    assign memory[5014] = 12'h890;
    assign memory[5015] = 12'hbb0;
    assign memory[5016] = 12'h780;
    assign memory[5017] = 12'h670;
    assign memory[5018] = 12'h890;
    assign memory[5019] = 12'h670;
    assign memory[5020] = 12'hbb0;
    assign memory[5021] = 12'hbb0;
    assign memory[5022] = 12'hbb0;
    assign memory[5023] = 12'hbb0;
    assign memory[5024] = 12'h890;
    assign memory[5025] = 12'hbb0;
    assign memory[5026] = 12'h890;
    assign memory[5027] = 12'hbb0;
    assign memory[5028] = 12'h670;
    assign memory[5029] = 12'hbb0;
    assign memory[5030] = 12'hbb0;
    assign memory[5031] = 12'h670;
    assign memory[5032] = 12'h890;
    assign memory[5033] = 12'hbb0;
    assign memory[5034] = 12'h890;
    assign memory[5035] = 12'hbb0;
    assign memory[5036] = 12'h890;
    assign memory[5037] = 12'hbb0;
    assign memory[5038] = 12'h670;
    assign memory[5039] = 12'hbb0;
    assign memory[5040] = 12'hbb0;
    assign memory[5041] = 12'hbb0;
    assign memory[5042] = 12'h670;
    assign memory[5043] = 12'hbb0;
    assign memory[5044] = 12'hbb0;
    assign memory[5045] = 12'h890;
    assign memory[5046] = 12'hbb0;
    assign memory[5047] = 12'hbb0;
    assign memory[5048] = 12'h780;
    assign memory[5049] = 12'h670;
    assign memory[5050] = 12'h890;
    assign memory[5051] = 12'hbb0;
    assign memory[5052] = 12'hbb0;
    assign memory[5053] = 12'hbb0;
    assign memory[5054] = 12'hbb0;
    assign memory[5055] = 12'hbb0;
    assign memory[5056] = 12'h890;
    assign memory[5057] = 12'hbb0;
    assign memory[5058] = 12'h890;
    assign memory[5059] = 12'hbb0;
    assign memory[5060] = 12'h670;
    assign memory[5061] = 12'hbb0;
    assign memory[5062] = 12'hbb0;
    assign memory[5063] = 12'h670;
    assign memory[5064] = 12'h890;
    assign memory[5065] = 12'hbb0;
    assign memory[5066] = 12'h890;
    assign memory[5067] = 12'hbb0;
    assign memory[5068] = 12'h890;
    assign memory[5069] = 12'h670;
    assign memory[5070] = 12'hbb0;
    assign memory[5071] = 12'hbb0;
    assign memory[5072] = 12'hbb0;
    assign memory[5073] = 12'hbb0;
    assign memory[5074] = 12'h670;
    assign memory[5075] = 12'hbb0;
    assign memory[5076] = 12'hbb0;
    assign memory[5077] = 12'h890;
    assign memory[5078] = 12'hbb0;
    assign memory[5079] = 12'hbb0;
    assign memory[5080] = 12'h780;
    assign memory[5081] = 12'h670;
    assign memory[5082] = 12'hbb0;
    assign memory[5083] = 12'hbb0;
    assign memory[5084] = 12'hbb0;
    assign memory[5085] = 12'hbb0;
    assign memory[5086] = 12'hbb0;
    assign memory[5087] = 12'hbb0;
    assign memory[5088] = 12'h890;
    assign memory[5089] = 12'hbb0;
    assign memory[5090] = 12'h890;
    assign memory[5091] = 12'hbb0;
    assign memory[5092] = 12'h670;
    assign memory[5093] = 12'hbb0;
    assign memory[5094] = 12'hbb0;
    assign memory[5095] = 12'hbb0;
    assign memory[5096] = 12'h890;
    assign memory[5097] = 12'hbb0;
    assign memory[5098] = 12'h890;
    assign memory[5099] = 12'hbb0;
    assign memory[5100] = 12'h890;
    assign memory[5101] = 12'h670;
    assign memory[5102] = 12'hbb0;
    assign memory[5103] = 12'hbb0;
    assign memory[5104] = 12'hbb0;
    assign memory[5105] = 12'hbb0;
    assign memory[5106] = 12'h670;
    assign memory[5107] = 12'hbb0;
    assign memory[5108] = 12'hbb0;
    assign memory[5109] = 12'h890;
    assign memory[5110] = 12'hbb0;
    assign memory[5111] = 12'hbb0;
    assign memory[5112] = 12'hbb0;
    assign memory[5113] = 12'h670;
    assign memory[5114] = 12'hbb0;
    assign memory[5115] = 12'hbb0;
    assign memory[5116] = 12'hbb0;
    assign memory[5117] = 12'hbb0;
    assign memory[5118] = 12'hbb0;
    assign memory[5119] = 12'hbb0;
    assign memory[5120] = 12'hd84;
    assign memory[5121] = 12'hd84;
    assign memory[5122] = 12'hd84;
    assign memory[5123] = 12'hd84;
    assign memory[5124] = 12'hd84;
    assign memory[5125] = 12'hd84;
    assign memory[5126] = 12'hd84;
    assign memory[5127] = 12'hd84;
    assign memory[5128] = 12'hd84;
    assign memory[5129] = 12'hd84;
    assign memory[5130] = 12'hd84;
    assign memory[5131] = 12'hd84;
    assign memory[5132] = 12'hd74;
    assign memory[5133] = 12'hd85;
    assign memory[5134] = 12'hd84;
    assign memory[5135] = 12'hd84;
    assign memory[5136] = 12'hd84;
    assign memory[5137] = 12'hd84;
    assign memory[5138] = 12'hd84;
    assign memory[5139] = 12'hd74;
    assign memory[5140] = 12'hd84;
    assign memory[5141] = 12'hd84;
    assign memory[5142] = 12'hd84;
    assign memory[5143] = 12'hd84;
    assign memory[5144] = 12'hd84;
    assign memory[5145] = 12'hd84;
    assign memory[5146] = 12'hd84;
    assign memory[5147] = 12'hd84;
    assign memory[5148] = 12'hd84;
    assign memory[5149] = 12'hd84;
    assign memory[5150] = 12'hd84;
    assign memory[5151] = 12'hd84;
    assign memory[5152] = 12'hd84;
    assign memory[5153] = 12'hd84;
    assign memory[5154] = 12'hd74;
    assign memory[5155] = 12'hd84;
    assign memory[5156] = 12'hc94;
    assign memory[5157] = 12'hd84;
    assign memory[5158] = 12'hd84;
    assign memory[5159] = 12'hd74;
    assign memory[5160] = 12'hd85;
    assign memory[5161] = 12'hc94;
    assign memory[5162] = 12'hd84;
    assign memory[5163] = 12'hd84;
    assign memory[5164] = 12'hd84;
    assign memory[5165] = 12'hd85;
    assign memory[5166] = 12'hd74;
    assign memory[5167] = 12'hd84;
    assign memory[5168] = 12'hd84;
    assign memory[5169] = 12'hd84;
    assign memory[5170] = 12'hc94;
    assign memory[5171] = 12'hd84;
    assign memory[5172] = 12'hd84;
    assign memory[5173] = 12'hc94;
    assign memory[5174] = 12'hd84;
    assign memory[5175] = 12'hc94;
    assign memory[5176] = 12'hd84;
    assign memory[5177] = 12'hc94;
    assign memory[5178] = 12'hd84;
    assign memory[5179] = 12'hd84;
    assign memory[5180] = 12'hd74;
    assign memory[5181] = 12'hd84;
    assign memory[5182] = 12'hd84;
    assign memory[5183] = 12'hd84;
    assign memory[5184] = 12'hd84;
    assign memory[5185] = 12'hd84;
    assign memory[5186] = 12'hd84;
    assign memory[5187] = 12'hd74;
    assign memory[5188] = 12'hd84;
    assign memory[5189] = 12'hd84;
    assign memory[5190] = 12'hd84;
    assign memory[5191] = 12'hd84;
    assign memory[5192] = 12'hd84;
    assign memory[5193] = 12'hd84;
    assign memory[5194] = 12'hd84;
    assign memory[5195] = 12'hd84;
    assign memory[5196] = 12'hd84;
    assign memory[5197] = 12'hd84;
    assign memory[5198] = 12'hd84;
    assign memory[5199] = 12'hc94;
    assign memory[5200] = 12'hd84;
    assign memory[5201] = 12'hd84;
    assign memory[5202] = 12'hd74;
    assign memory[5203] = 12'hd74;
    assign memory[5204] = 12'hd84;
    assign memory[5205] = 12'hd84;
    assign memory[5206] = 12'hd85;
    assign memory[5207] = 12'hd84;
    assign memory[5208] = 12'hc94;
    assign memory[5209] = 12'hd84;
    assign memory[5210] = 12'hd84;
    assign memory[5211] = 12'hd84;
    assign memory[5212] = 12'hd84;
    assign memory[5213] = 12'hd84;
    assign memory[5214] = 12'hd84;
    assign memory[5215] = 12'hd84;
    assign memory[5216] = 12'hd84;
    assign memory[5217] = 12'hd84;
    assign memory[5218] = 12'hc94;
    assign memory[5219] = 12'hc94;
    assign memory[5220] = 12'hd74;
    assign memory[5221] = 12'hd84;
    assign memory[5222] = 12'hd84;
    assign memory[5223] = 12'hd84;
    assign memory[5224] = 12'hd84;
    assign memory[5225] = 12'hd84;
    assign memory[5226] = 12'hd84;
    assign memory[5227] = 12'hd84;
    assign memory[5228] = 12'hc94;
    assign memory[5229] = 12'hd84;
    assign memory[5230] = 12'hd84;
    assign memory[5231] = 12'hd74;
    assign memory[5232] = 12'hd84;
    assign memory[5233] = 12'hc94;
    assign memory[5234] = 12'hd85;
    assign memory[5235] = 12'hd74;
    assign memory[5236] = 12'hd84;
    assign memory[5237] = 12'hd84;
    assign memory[5238] = 12'hd84;
    assign memory[5239] = 12'hd84;
    assign memory[5240] = 12'hd84;
    assign memory[5241] = 12'hd84;
    assign memory[5242] = 12'hd84;
    assign memory[5243] = 12'hd84;
    assign memory[5244] = 12'hd84;
    assign memory[5245] = 12'hd84;
    assign memory[5246] = 12'hd85;
    assign memory[5247] = 12'hd84;
    assign memory[5248] = 12'hd84;
    assign memory[5249] = 12'hd84;
    assign memory[5250] = 12'hd84;
    assign memory[5251] = 12'hc94;
    assign memory[5252] = 12'hd84;
    assign memory[5253] = 12'hc94;
    assign memory[5254] = 12'hd84;
    assign memory[5255] = 12'hd84;
    assign memory[5256] = 12'hd84;
    assign memory[5257] = 12'hd84;
    assign memory[5258] = 12'hd84;
    assign memory[5259] = 12'hd84;
    assign memory[5260] = 12'hd84;
    assign memory[5261] = 12'hd84;
    assign memory[5262] = 12'hd84;
    assign memory[5263] = 12'hd84;
    assign memory[5264] = 12'hd84;
    assign memory[5265] = 12'hd84;
    assign memory[5266] = 12'hd84;
    assign memory[5267] = 12'hd84;
    assign memory[5268] = 12'hd84;
    assign memory[5269] = 12'hd84;
    assign memory[5270] = 12'hc94;
    assign memory[5271] = 12'hd74;
    assign memory[5272] = 12'hd84;
    assign memory[5273] = 12'hd84;
    assign memory[5274] = 12'hd84;
    assign memory[5275] = 12'hd84;
    assign memory[5276] = 12'hd84;
    assign memory[5277] = 12'hd84;
    assign memory[5278] = 12'hd84;
    assign memory[5279] = 12'hd84;
    assign memory[5280] = 12'hd84;
    assign memory[5281] = 12'hc94;
    assign memory[5282] = 12'hd84;
    assign memory[5283] = 12'hc94;
    assign memory[5284] = 12'hd84;
    assign memory[5285] = 12'hd84;
    assign memory[5286] = 12'hd84;
    assign memory[5287] = 12'hd84;
    assign memory[5288] = 12'hd84;
    assign memory[5289] = 12'hd84;
    assign memory[5290] = 12'hc94;
    assign memory[5291] = 12'hd84;
    assign memory[5292] = 12'hd84;
    assign memory[5293] = 12'hd84;
    assign memory[5294] = 12'hd84;
    assign memory[5295] = 12'hd84;
    assign memory[5296] = 12'hc94;
    assign memory[5297] = 12'hd84;
    assign memory[5298] = 12'hd74;
    assign memory[5299] = 12'hd84;
    assign memory[5300] = 12'hd84;
    assign memory[5301] = 12'hc94;
    assign memory[5302] = 12'hd84;
    assign memory[5303] = 12'hd74;
    assign memory[5304] = 12'hd84;
    assign memory[5305] = 12'hd84;
    assign memory[5306] = 12'hd84;
    assign memory[5307] = 12'hd84;
    assign memory[5308] = 12'hd84;
    assign memory[5309] = 12'hd84;
    assign memory[5310] = 12'hd84;
    assign memory[5311] = 12'hd84;
    assign memory[5312] = 12'hd84;
    assign memory[5313] = 12'hd84;
    assign memory[5314] = 12'hd84;
    assign memory[5315] = 12'hd84;
    assign memory[5316] = 12'hd74;
    assign memory[5317] = 12'hd84;
    assign memory[5318] = 12'hd84;
    assign memory[5319] = 12'hd84;
    assign memory[5320] = 12'hd84;
    assign memory[5321] = 12'hd84;
    assign memory[5322] = 12'hd84;
    assign memory[5323] = 12'hd84;
    assign memory[5324] = 12'hd85;
    assign memory[5325] = 12'hd74;
    assign memory[5326] = 12'hd84;
    assign memory[5327] = 12'hd84;
    assign memory[5328] = 12'hd84;
    assign memory[5329] = 12'hd84;
    assign memory[5330] = 12'hd84;
    assign memory[5331] = 12'hc94;
    assign memory[5332] = 12'hd84;
    assign memory[5333] = 12'hccc;
    assign memory[5334] = 12'haaa;
    assign memory[5335] = 12'hd84;
    assign memory[5336] = 12'hd84;
    assign memory[5337] = 12'hd84;
    assign memory[5338] = 12'hd84;
    assign memory[5339] = 12'hd74;
    assign memory[5340] = 12'hd84;
    assign memory[5341] = 12'hd84;
    assign memory[5342] = 12'hd84;
    assign memory[5343] = 12'hd84;
    assign memory[5344] = 12'hd84;
    assign memory[5345] = 12'hd84;
    assign memory[5346] = 12'hd84;
    assign memory[5347] = 12'hd84;
    assign memory[5348] = 12'hc94;
    assign memory[5349] = 12'hd84;
    assign memory[5350] = 12'hd84;
    assign memory[5351] = 12'hd84;
    assign memory[5352] = 12'hd84;
    assign memory[5353] = 12'hd85;
    assign memory[5354] = 12'hd84;
    assign memory[5355] = 12'hc94;
    assign memory[5356] = 12'hd74;
    assign memory[5357] = 12'hd84;
    assign memory[5358] = 12'hd84;
    assign memory[5359] = 12'hd84;
    assign memory[5360] = 12'hc94;
    assign memory[5361] = 12'hd84;
    assign memory[5362] = 12'hd74;
    assign memory[5363] = 12'hd84;
    assign memory[5364] = 12'hccc;
    assign memory[5365] = 12'hccc;
    assign memory[5366] = 12'hccc;
    assign memory[5367] = 12'haaa;
    assign memory[5368] = 12'hc94;
    assign memory[5369] = 12'hd84;
    assign memory[5370] = 12'hd84;
    assign memory[5371] = 12'hd84;
    assign memory[5372] = 12'hd84;
    assign memory[5373] = 12'hd84;
    assign memory[5374] = 12'hd84;
    assign memory[5375] = 12'hd84;
    assign memory[5376] = 12'hd84;
    assign memory[5377] = 12'hd84;
    assign memory[5378] = 12'hd84;
    assign memory[5379] = 12'hd85;
    assign memory[5380] = 12'hd84;
    assign memory[5381] = 12'hd84;
    assign memory[5382] = 12'hd84;
    assign memory[5383] = 12'hd84;
    assign memory[5384] = 12'hd84;
    assign memory[5385] = 12'hd84;
    assign memory[5386] = 12'hd85;
    assign memory[5387] = 12'hd74;
    assign memory[5388] = 12'hd84;
    assign memory[5389] = 12'hd84;
    assign memory[5390] = 12'hd84;
    assign memory[5391] = 12'hc94;
    assign memory[5392] = 12'hc94;
    assign memory[5393] = 12'hd84;
    assign memory[5394] = 12'hd84;
    assign memory[5395] = 12'hd84;
    assign memory[5396] = 12'hccc;
    assign memory[5397] = 12'hccc;
    assign memory[5398] = 12'hccc;
    assign memory[5399] = 12'haaa;
    assign memory[5400] = 12'haaa;
    assign memory[5401] = 12'hc94;
    assign memory[5402] = 12'hd84;
    assign memory[5403] = 12'hd84;
    assign memory[5404] = 12'hd84;
    assign memory[5405] = 12'hd84;
    assign memory[5406] = 12'hd84;
    assign memory[5407] = 12'hd84;
    assign memory[5408] = 12'hd84;
    assign memory[5409] = 12'hc94;
    assign memory[5410] = 12'hd84;
    assign memory[5411] = 12'hd74;
    assign memory[5412] = 12'hd84;
    assign memory[5413] = 12'hd84;
    assign memory[5414] = 12'hd84;
    assign memory[5415] = 12'hd84;
    assign memory[5416] = 12'hd84;
    assign memory[5417] = 12'hd84;
    assign memory[5418] = 12'hd84;
    assign memory[5419] = 12'hd74;
    assign memory[5420] = 12'hd84;
    assign memory[5421] = 12'hd85;
    assign memory[5422] = 12'hd84;
    assign memory[5423] = 12'hd84;
    assign memory[5424] = 12'hbe1;
    assign memory[5425] = 12'hd84;
    assign memory[5426] = 12'hd84;
    assign memory[5427] = 12'hccc;
    assign memory[5428] = 12'hccc;
    assign memory[5429] = 12'hccc;
    assign memory[5430] = 12'hccc;
    assign memory[5431] = 12'haaa;
    assign memory[5432] = 12'haaa;
    assign memory[5433] = 12'hd84;
    assign memory[5434] = 12'hd84;
    assign memory[5435] = 12'hd84;
    assign memory[5436] = 12'hd74;
    assign memory[5437] = 12'hd84;
    assign memory[5438] = 12'hd84;
    assign memory[5439] = 12'hd74;
    assign memory[5440] = 12'hd84;
    assign memory[5441] = 12'hd84;
    assign memory[5442] = 12'hd84;
    assign memory[5443] = 12'hd84;
    assign memory[5444] = 12'hd84;
    assign memory[5445] = 12'hd84;
    assign memory[5446] = 12'hd84;
    assign memory[5447] = 12'hd84;
    assign memory[5448] = 12'hd84;
    assign memory[5449] = 12'hd84;
    assign memory[5450] = 12'hd84;
    assign memory[5451] = 12'hc94;
    assign memory[5452] = 12'hd84;
    assign memory[5453] = 12'hd84;
    assign memory[5454] = 12'hd84;
    assign memory[5455] = 12'hd84;
    assign memory[5456] = 12'hbe1;
    assign memory[5457] = 12'hbe1;
    assign memory[5458] = 12'hd84;
    assign memory[5459] = 12'hbe1;
    assign memory[5460] = 12'hbe1;
    assign memory[5461] = 12'hbe1;
    assign memory[5462] = 12'hd84;
    assign memory[5463] = 12'hd74;
    assign memory[5464] = 12'hd74;
    assign memory[5465] = 12'hd85;
    assign memory[5466] = 12'hd84;
    assign memory[5467] = 12'hd84;
    assign memory[5468] = 12'hd84;
    assign memory[5469] = 12'hd84;
    assign memory[5470] = 12'hd85;
    assign memory[5471] = 12'hd84;
    assign memory[5472] = 12'hd84;
    assign memory[5473] = 12'hd84;
    assign memory[5474] = 12'hd84;
    assign memory[5475] = 12'hc94;
    assign memory[5476] = 12'hd85;
    assign memory[5477] = 12'hd84;
    assign memory[5478] = 12'hd84;
    assign memory[5479] = 12'hd84;
    assign memory[5480] = 12'hc94;
    assign memory[5481] = 12'hc94;
    assign memory[5482] = 12'hd84;
    assign memory[5483] = 12'hd84;
    assign memory[5484] = 12'hd84;
    assign memory[5485] = 12'hd84;
    assign memory[5486] = 12'hd84;
    assign memory[5487] = 12'hc94;
    assign memory[5488] = 12'hbe1;
    assign memory[5489] = 12'hbe1;
    assign memory[5490] = 12'hbe1;
    assign memory[5491] = 12'hbe1;
    assign memory[5492] = 12'hbe1;
    assign memory[5493] = 12'hbe1;
    assign memory[5494] = 12'hd85;
    assign memory[5495] = 12'hd84;
    assign memory[5496] = 12'hd85;
    assign memory[5497] = 12'hc94;
    assign memory[5498] = 12'hc94;
    assign memory[5499] = 12'hd84;
    assign memory[5500] = 12'hd74;
    assign memory[5501] = 12'hd84;
    assign memory[5502] = 12'hc94;
    assign memory[5503] = 12'hd84;
    assign memory[5504] = 12'hc94;
    assign memory[5505] = 12'hc94;
    assign memory[5506] = 12'hd84;
    assign memory[5507] = 12'hd84;
    assign memory[5508] = 12'hd85;
    assign memory[5509] = 12'hd85;
    assign memory[5510] = 12'hd85;
    assign memory[5511] = 12'hd84;
    assign memory[5512] = 12'hd84;
    assign memory[5513] = 12'hd84;
    assign memory[5514] = 12'hd74;
    assign memory[5515] = 12'hd84;
    assign memory[5516] = 12'hd84;
    assign memory[5517] = 12'hd84;
    assign memory[5518] = 12'hd84;
    assign memory[5519] = 12'hd84;
    assign memory[5520] = 12'hc94;
    assign memory[5521] = 12'hc94;
    assign memory[5522] = 12'hd84;
    assign memory[5523] = 12'hc94;
    assign memory[5524] = 12'hd84;
    assign memory[5525] = 12'hc94;
    assign memory[5526] = 12'hc94;
    assign memory[5527] = 12'hd84;
    assign memory[5528] = 12'hd84;
    assign memory[5529] = 12'hd84;
    assign memory[5530] = 12'hd84;
    assign memory[5531] = 12'hd74;
    assign memory[5532] = 12'hd74;
    assign memory[5533] = 12'hd84;
    assign memory[5534] = 12'hd84;
    assign memory[5535] = 12'hd84;
    assign memory[5536] = 12'hd84;
    assign memory[5537] = 12'hd84;
    assign memory[5538] = 12'hd84;
    assign memory[5539] = 12'hd84;
    assign memory[5540] = 12'hd84;
    assign memory[5541] = 12'hd84;
    assign memory[5542] = 12'hc94;
    assign memory[5543] = 12'hc94;
    assign memory[5544] = 12'hd84;
    assign memory[5545] = 12'hd84;
    assign memory[5546] = 12'hd84;
    assign memory[5547] = 12'hd84;
    assign memory[5548] = 12'hd84;
    assign memory[5549] = 12'hd84;
    assign memory[5550] = 12'hd85;
    assign memory[5551] = 12'hd84;
    assign memory[5552] = 12'hc94;
    assign memory[5553] = 12'hc94;
    assign memory[5554] = 12'hd84;
    assign memory[5555] = 12'hc94;
    assign memory[5556] = 12'hd84;
    assign memory[5557] = 12'hc94;
    assign memory[5558] = 12'hc94;
    assign memory[5559] = 12'hd84;
    assign memory[5560] = 12'hd84;
    assign memory[5561] = 12'hd84;
    assign memory[5562] = 12'hd84;
    assign memory[5563] = 12'hd84;
    assign memory[5564] = 12'hd84;
    assign memory[5565] = 12'hd84;
    assign memory[5566] = 12'hd84;
    assign memory[5567] = 12'hd74;
    assign memory[5568] = 12'hd84;
    assign memory[5569] = 12'hd84;
    assign memory[5570] = 12'hd84;
    assign memory[5571] = 12'hd84;
    assign memory[5572] = 12'hd84;
    assign memory[5573] = 12'hd84;
    assign memory[5574] = 12'hd84;
    assign memory[5575] = 12'hd84;
    assign memory[5576] = 12'hd84;
    assign memory[5577] = 12'hd84;
    assign memory[5578] = 12'hd84;
    assign memory[5579] = 12'hd84;
    assign memory[5580] = 12'hd84;
    assign memory[5581] = 12'hd84;
    assign memory[5582] = 12'hd84;
    assign memory[5583] = 12'hd74;
    assign memory[5584] = 12'hc94;
    assign memory[5585] = 12'hd84;
    assign memory[5586] = 12'hd84;
    assign memory[5587] = 12'hc94;
    assign memory[5588] = 12'hd84;
    assign memory[5589] = 12'hd84;
    assign memory[5590] = 12'hd84;
    assign memory[5591] = 12'hd74;
    assign memory[5592] = 12'hd84;
    assign memory[5593] = 12'hd84;
    assign memory[5594] = 12'hd74;
    assign memory[5595] = 12'hd84;
    assign memory[5596] = 12'hd84;
    assign memory[5597] = 12'hd84;
    assign memory[5598] = 12'hd84;
    assign memory[5599] = 12'hd84;
    assign memory[5600] = 12'hd84;
    assign memory[5601] = 12'hd84;
    assign memory[5602] = 12'hd84;
    assign memory[5603] = 12'hd84;
    assign memory[5604] = 12'hd84;
    assign memory[5605] = 12'hd84;
    assign memory[5606] = 12'hc94;
    assign memory[5607] = 12'hd84;
    assign memory[5608] = 12'hd84;
    assign memory[5609] = 12'hd84;
    assign memory[5610] = 12'hd84;
    assign memory[5611] = 12'hd84;
    assign memory[5612] = 12'hd84;
    assign memory[5613] = 12'hd85;
    assign memory[5614] = 12'hd84;
    assign memory[5615] = 12'hd84;
    assign memory[5616] = 12'hd84;
    assign memory[5617] = 12'hd84;
    assign memory[5618] = 12'hd85;
    assign memory[5619] = 12'hd84;
    assign memory[5620] = 12'hd84;
    assign memory[5621] = 12'hd84;
    assign memory[5622] = 12'hd84;
    assign memory[5623] = 12'hc94;
    assign memory[5624] = 12'hd74;
    assign memory[5625] = 12'hd84;
    assign memory[5626] = 12'hc94;
    assign memory[5627] = 12'hd84;
    assign memory[5628] = 12'hd84;
    assign memory[5629] = 12'hd84;
    assign memory[5630] = 12'hd74;
    assign memory[5631] = 12'hd84;
    assign memory[5632] = 12'hd84;
    assign memory[5633] = 12'hd84;
    assign memory[5634] = 12'hd84;
    assign memory[5635] = 12'hd84;
    assign memory[5636] = 12'hd84;
    assign memory[5637] = 12'hc94;
    assign memory[5638] = 12'hd84;
    assign memory[5639] = 12'hd84;
    assign memory[5640] = 12'hd74;
    assign memory[5641] = 12'hd84;
    assign memory[5642] = 12'hd74;
    assign memory[5643] = 12'hd84;
    assign memory[5644] = 12'hd84;
    assign memory[5645] = 12'hd74;
    assign memory[5646] = 12'hd84;
    assign memory[5647] = 12'hd84;
    assign memory[5648] = 12'hd84;
    assign memory[5649] = 12'hd84;
    assign memory[5650] = 12'hd84;
    assign memory[5651] = 12'hd84;
    assign memory[5652] = 12'hd84;
    assign memory[5653] = 12'hd84;
    assign memory[5654] = 12'hd84;
    assign memory[5655] = 12'hd74;
    assign memory[5656] = 12'hc94;
    assign memory[5657] = 12'hd84;
    assign memory[5658] = 12'hd84;
    assign memory[5659] = 12'hd85;
    assign memory[5660] = 12'hd84;
    assign memory[5661] = 12'hd84;
    assign memory[5662] = 12'hd84;
    assign memory[5663] = 12'hc94;
    assign memory[5664] = 12'hd74;
    assign memory[5665] = 12'hd84;
    assign memory[5666] = 12'hd84;
    assign memory[5667] = 12'hd84;
    assign memory[5668] = 12'hd84;
    assign memory[5669] = 12'hd84;
    assign memory[5670] = 12'hd84;
    assign memory[5671] = 12'hd84;
    assign memory[5672] = 12'hd84;
    assign memory[5673] = 12'hd84;
    assign memory[5674] = 12'hd84;
    assign memory[5675] = 12'hd74;
    assign memory[5676] = 12'hd84;
    assign memory[5677] = 12'hd84;
    assign memory[5678] = 12'hd74;
    assign memory[5679] = 12'hd84;
    assign memory[5680] = 12'hd84;
    assign memory[5681] = 12'hd74;
    assign memory[5682] = 12'hd74;
    assign memory[5683] = 12'hd74;
    assign memory[5684] = 12'hd84;
    assign memory[5685] = 12'hd84;
    assign memory[5686] = 12'hd84;
    assign memory[5687] = 12'hd84;
    assign memory[5688] = 12'hd74;
    assign memory[5689] = 12'hd84;
    assign memory[5690] = 12'hd84;
    assign memory[5691] = 12'hd84;
    assign memory[5692] = 12'hd84;
    assign memory[5693] = 12'hd84;
    assign memory[5694] = 12'hd84;
    assign memory[5695] = 12'hd84;
    assign memory[5696] = 12'hd84;
    assign memory[5697] = 12'hd84;
    assign memory[5698] = 12'hd84;
    assign memory[5699] = 12'hd84;
    assign memory[5700] = 12'hd84;
    assign memory[5701] = 12'hd84;
    assign memory[5702] = 12'hd74;
    assign memory[5703] = 12'hd84;
    assign memory[5704] = 12'hd84;
    assign memory[5705] = 12'hd84;
    assign memory[5706] = 12'hd84;
    assign memory[5707] = 12'hd84;
    assign memory[5708] = 12'hd84;
    assign memory[5709] = 12'hd84;
    assign memory[5710] = 12'hd84;
    assign memory[5711] = 12'hd84;
    assign memory[5712] = 12'hd84;
    assign memory[5713] = 12'hd84;
    assign memory[5714] = 12'hd84;
    assign memory[5715] = 12'hc94;
    assign memory[5716] = 12'hd84;
    assign memory[5717] = 12'hd84;
    assign memory[5718] = 12'hd84;
    assign memory[5719] = 12'hd74;
    assign memory[5720] = 12'hc94;
    assign memory[5721] = 12'hd84;
    assign memory[5722] = 12'hd84;
    assign memory[5723] = 12'hd84;
    assign memory[5724] = 12'hd84;
    assign memory[5725] = 12'hd84;
    assign memory[5726] = 12'hc94;
    assign memory[5727] = 12'hd84;
    assign memory[5728] = 12'hc94;
    assign memory[5729] = 12'hc94;
    assign memory[5730] = 12'hd84;
    assign memory[5731] = 12'hd84;
    assign memory[5732] = 12'hd84;
    assign memory[5733] = 12'hd84;
    assign memory[5734] = 12'hd84;
    assign memory[5735] = 12'hd84;
    assign memory[5736] = 12'hd84;
    assign memory[5737] = 12'hd84;
    assign memory[5738] = 12'hd84;
    assign memory[5739] = 12'hd84;
    assign memory[5740] = 12'hd74;
    assign memory[5741] = 12'hc94;
    assign memory[5742] = 12'hd84;
    assign memory[5743] = 12'hd84;
    assign memory[5744] = 12'hd74;
    assign memory[5745] = 12'hd84;
    assign memory[5746] = 12'hd74;
    assign memory[5747] = 12'hd84;
    assign memory[5748] = 12'hd84;
    assign memory[5749] = 12'hc94;
    assign memory[5750] = 12'hd84;
    assign memory[5751] = 12'hc94;
    assign memory[5752] = 12'hd84;
    assign memory[5753] = 12'hd84;
    assign memory[5754] = 12'hd84;
    assign memory[5755] = 12'hc94;
    assign memory[5756] = 12'hd84;
    assign memory[5757] = 12'hd84;
    assign memory[5758] = 12'hd84;
    assign memory[5759] = 12'hd84;
    assign memory[5760] = 12'hd84;
    assign memory[5761] = 12'hd84;
    assign memory[5762] = 12'hd84;
    assign memory[5763] = 12'hd84;
    assign memory[5764] = 12'hd84;
    assign memory[5765] = 12'hd84;
    assign memory[5766] = 12'hd84;
    assign memory[5767] = 12'hd84;
    assign memory[5768] = 12'hd84;
    assign memory[5769] = 12'hd84;
    assign memory[5770] = 12'hd84;
    assign memory[5771] = 12'hd84;
    assign memory[5772] = 12'hd84;
    assign memory[5773] = 12'hd84;
    assign memory[5774] = 12'hd84;
    assign memory[5775] = 12'hd84;
    assign memory[5776] = 12'hc94;
    assign memory[5777] = 12'hd84;
    assign memory[5778] = 12'hd84;
    assign memory[5779] = 12'hd84;
    assign memory[5780] = 12'hd84;
    assign memory[5781] = 12'hd84;
    assign memory[5782] = 12'hd84;
    assign memory[5783] = 12'hd84;
    assign memory[5784] = 12'hd84;
    assign memory[5785] = 12'hd84;
    assign memory[5786] = 12'hd84;
    assign memory[5787] = 12'hd84;
    assign memory[5788] = 12'hd84;
    assign memory[5789] = 12'hd84;
    assign memory[5790] = 12'hd84;
    assign memory[5791] = 12'hd84;
    assign memory[5792] = 12'hc94;
    assign memory[5793] = 12'hd84;
    assign memory[5794] = 12'hd84;
    assign memory[5795] = 12'hd84;
    assign memory[5796] = 12'hd84;
    assign memory[5797] = 12'hd84;
    assign memory[5798] = 12'hd84;
    assign memory[5799] = 12'hccc;
    assign memory[5800] = 12'haaa;
    assign memory[5801] = 12'hd84;
    assign memory[5802] = 12'hd84;
    assign memory[5803] = 12'hd84;
    assign memory[5804] = 12'hd84;
    assign memory[5805] = 12'hd84;
    assign memory[5806] = 12'hd84;
    assign memory[5807] = 12'hd84;
    assign memory[5808] = 12'hd84;
    assign memory[5809] = 12'hd84;
    assign memory[5810] = 12'hd84;
    assign memory[5811] = 12'hd84;
    assign memory[5812] = 12'hd84;
    assign memory[5813] = 12'hd84;
    assign memory[5814] = 12'hd84;
    assign memory[5815] = 12'hd84;
    assign memory[5816] = 12'hd84;
    assign memory[5817] = 12'hd84;
    assign memory[5818] = 12'hd84;
    assign memory[5819] = 12'hd84;
    assign memory[5820] = 12'hd84;
    assign memory[5821] = 12'hd84;
    assign memory[5822] = 12'hd84;
    assign memory[5823] = 12'hd84;
    assign memory[5824] = 12'hd84;
    assign memory[5825] = 12'hd84;
    assign memory[5826] = 12'hd84;
    assign memory[5827] = 12'hd84;
    assign memory[5828] = 12'hd84;
    assign memory[5829] = 12'hd84;
    assign memory[5830] = 12'hccc;
    assign memory[5831] = 12'hccc;
    assign memory[5832] = 12'haaa;
    assign memory[5833] = 12'haaa;
    assign memory[5834] = 12'hd74;
    assign memory[5835] = 12'hd84;
    assign memory[5836] = 12'hd84;
    assign memory[5837] = 12'hd84;
    assign memory[5838] = 12'hd84;
    assign memory[5839] = 12'hd84;
    assign memory[5840] = 12'hc94;
    assign memory[5841] = 12'hd84;
    assign memory[5842] = 12'hd84;
    assign memory[5843] = 12'hd74;
    assign memory[5844] = 12'hd84;
    assign memory[5845] = 12'hd84;
    assign memory[5846] = 12'hd84;
    assign memory[5847] = 12'hd84;
    assign memory[5848] = 12'hd84;
    assign memory[5849] = 12'hd84;
    assign memory[5850] = 12'hd84;
    assign memory[5851] = 12'hd84;
    assign memory[5852] = 12'hd84;
    assign memory[5853] = 12'hd84;
    assign memory[5854] = 12'hd84;
    assign memory[5855] = 12'hd84;
    assign memory[5856] = 12'hd84;
    assign memory[5857] = 12'hd84;
    assign memory[5858] = 12'hd84;
    assign memory[5859] = 12'hd84;
    assign memory[5860] = 12'hd84;
    assign memory[5861] = 12'hccc;
    assign memory[5862] = 12'hccc;
    assign memory[5863] = 12'hccc;
    assign memory[5864] = 12'hccc;
    assign memory[5865] = 12'haaa;
    assign memory[5866] = 12'haaa;
    assign memory[5867] = 12'hc94;
    assign memory[5868] = 12'hd84;
    assign memory[5869] = 12'hd84;
    assign memory[5870] = 12'hd84;
    assign memory[5871] = 12'hbe1;
    assign memory[5872] = 12'hd84;
    assign memory[5873] = 12'hbe1;
    assign memory[5874] = 12'hd84;
    assign memory[5875] = 12'hd84;
    assign memory[5876] = 12'hd84;
    assign memory[5877] = 12'hd84;
    assign memory[5878] = 12'hd84;
    assign memory[5879] = 12'hd84;
    assign memory[5880] = 12'hd84;
    assign memory[5881] = 12'hd84;
    assign memory[5882] = 12'hd84;
    assign memory[5883] = 12'hd84;
    assign memory[5884] = 12'hd84;
    assign memory[5885] = 12'hd84;
    assign memory[5886] = 12'hd84;
    assign memory[5887] = 12'hd84;
    assign memory[5888] = 12'hd84;
    assign memory[5889] = 12'hd84;
    assign memory[5890] = 12'hd84;
    assign memory[5891] = 12'hd84;
    assign memory[5892] = 12'hd74;
    assign memory[5893] = 12'hccc;
    assign memory[5894] = 12'hccc;
    assign memory[5895] = 12'hccc;
    assign memory[5896] = 12'hccc;
    assign memory[5897] = 12'haaa;
    assign memory[5898] = 12'hd74;
    assign memory[5899] = 12'hd84;
    assign memory[5900] = 12'hd84;
    assign memory[5901] = 12'hbe1;
    assign memory[5902] = 12'hbe1;
    assign memory[5903] = 12'hbe1;
    assign memory[5904] = 12'hbe1;
    assign memory[5905] = 12'hbe1;
    assign memory[5906] = 12'hbe1;
    assign memory[5907] = 12'hd84;
    assign memory[5908] = 12'hd84;
    assign memory[5909] = 12'hd84;
    assign memory[5910] = 12'hd74;
    assign memory[5911] = 12'hd84;
    assign memory[5912] = 12'hd84;
    assign memory[5913] = 12'hd84;
    assign memory[5914] = 12'hd84;
    assign memory[5915] = 12'hc94;
    assign memory[5916] = 12'hd84;
    assign memory[5917] = 12'hd84;
    assign memory[5918] = 12'hd84;
    assign memory[5919] = 12'hd84;
    assign memory[5920] = 12'hd84;
    assign memory[5921] = 12'hd84;
    assign memory[5922] = 12'hd84;
    assign memory[5923] = 12'hd84;
    assign memory[5924] = 12'hd84;
    assign memory[5925] = 12'hd84;
    assign memory[5926] = 12'hd85;
    assign memory[5927] = 12'hc94;
    assign memory[5928] = 12'hd84;
    assign memory[5929] = 12'hd84;
    assign memory[5930] = 12'hd74;
    assign memory[5931] = 12'hd74;
    assign memory[5932] = 12'hd85;
    assign memory[5933] = 12'hd84;
    assign memory[5934] = 12'hc94;
    assign memory[5935] = 12'hc94;
    assign memory[5936] = 12'hd84;
    assign memory[5937] = 12'hd84;
    assign memory[5938] = 12'hd84;
    assign memory[5939] = 12'hd84;
    assign memory[5940] = 12'hd74;
    assign memory[5941] = 12'hd85;
    assign memory[5942] = 12'hd84;
    assign memory[5943] = 12'hd84;
    assign memory[5944] = 12'hd84;
    assign memory[5945] = 12'hd84;
    assign memory[5946] = 12'hd84;
    assign memory[5947] = 12'hd84;
    assign memory[5948] = 12'hd84;
    assign memory[5949] = 12'hd84;
    assign memory[5950] = 12'hd84;
    assign memory[5951] = 12'hd84;
    assign memory[5952] = 12'hd84;
    assign memory[5953] = 12'hd84;
    assign memory[5954] = 12'hd84;
    assign memory[5955] = 12'hc94;
    assign memory[5956] = 12'hd74;
    assign memory[5957] = 12'hd84;
    assign memory[5958] = 12'hd84;
    assign memory[5959] = 12'hc94;
    assign memory[5960] = 12'hd84;
    assign memory[5961] = 12'hd84;
    assign memory[5962] = 12'hd84;
    assign memory[5963] = 12'hd84;
    assign memory[5964] = 12'hd84;
    assign memory[5965] = 12'hd84;
    assign memory[5966] = 12'hd84;
    assign memory[5967] = 12'hd84;
    assign memory[5968] = 12'hd84;
    assign memory[5969] = 12'hd84;
    assign memory[5970] = 12'hc94;
    assign memory[5971] = 12'hd84;
    assign memory[5972] = 12'hc94;
    assign memory[5973] = 12'hd84;
    assign memory[5974] = 12'hd84;
    assign memory[5975] = 12'hd84;
    assign memory[5976] = 12'hd84;
    assign memory[5977] = 12'hd84;
    assign memory[5978] = 12'hd84;
    assign memory[5979] = 12'hd74;
    assign memory[5980] = 12'hd84;
    assign memory[5981] = 12'hd84;
    assign memory[5982] = 12'hd84;
    assign memory[5983] = 12'hd84;
    assign memory[5984] = 12'hd84;
    assign memory[5985] = 12'hd84;
    assign memory[5986] = 12'hd84;
    assign memory[5987] = 12'hd84;
    assign memory[5988] = 12'hd84;
    assign memory[5989] = 12'hd85;
    assign memory[5990] = 12'hd84;
    assign memory[5991] = 12'hd84;
    assign memory[5992] = 12'hd84;
    assign memory[5993] = 12'hd85;
    assign memory[5994] = 12'hd84;
    assign memory[5995] = 12'hd84;
    assign memory[5996] = 12'hc94;
    assign memory[5997] = 12'hc94;
    assign memory[5998] = 12'hd84;
    assign memory[5999] = 12'hd84;
    assign memory[6000] = 12'hd84;
    assign memory[6001] = 12'hd84;
    assign memory[6002] = 12'hd84;
    assign memory[6003] = 12'hd84;
    assign memory[6004] = 12'hd84;
    assign memory[6005] = 12'hd74;
    assign memory[6006] = 12'hd84;
    assign memory[6007] = 12'hd84;
    assign memory[6008] = 12'hd84;
    assign memory[6009] = 12'hd84;
    assign memory[6010] = 12'hd84;
    assign memory[6011] = 12'hd84;
    assign memory[6012] = 12'hc94;
    assign memory[6013] = 12'hd84;
    assign memory[6014] = 12'hd85;
    assign memory[6015] = 12'hd84;
    assign memory[6016] = 12'hd84;
    assign memory[6017] = 12'hc94;
    assign memory[6018] = 12'hd84;
    assign memory[6019] = 12'hc94;
    assign memory[6020] = 12'hd84;
    assign memory[6021] = 12'hd84;
    assign memory[6022] = 12'hd84;
    assign memory[6023] = 12'hd84;
    assign memory[6024] = 12'hd84;
    assign memory[6025] = 12'hd84;
    assign memory[6026] = 12'hd84;
    assign memory[6027] = 12'hd85;
    assign memory[6028] = 12'hd85;
    assign memory[6029] = 12'hd84;
    assign memory[6030] = 12'hd84;
    assign memory[6031] = 12'hd84;
    assign memory[6032] = 12'hd84;
    assign memory[6033] = 12'hc94;
    assign memory[6034] = 12'hd84;
    assign memory[6035] = 12'hd84;
    assign memory[6036] = 12'hd84;
    assign memory[6037] = 12'hd84;
    assign memory[6038] = 12'hd84;
    assign memory[6039] = 12'hd84;
    assign memory[6040] = 12'hd84;
    assign memory[6041] = 12'hd84;
    assign memory[6042] = 12'hd84;
    assign memory[6043] = 12'hd84;
    assign memory[6044] = 12'hd84;
    assign memory[6045] = 12'hd84;
    assign memory[6046] = 12'hd84;
    assign memory[6047] = 12'hd74;
    assign memory[6048] = 12'hd84;
    assign memory[6049] = 12'hd84;
    assign memory[6050] = 12'hd84;
    assign memory[6051] = 12'hd84;
    assign memory[6052] = 12'hd84;
    assign memory[6053] = 12'hd84;
    assign memory[6054] = 12'hd74;
    assign memory[6055] = 12'hd84;
    assign memory[6056] = 12'hc94;
    assign memory[6057] = 12'hd84;
    assign memory[6058] = 12'hd84;
    assign memory[6059] = 12'hd84;
    assign memory[6060] = 12'hd84;
    assign memory[6061] = 12'hd84;
    assign memory[6062] = 12'hd84;
    assign memory[6063] = 12'hd84;
    assign memory[6064] = 12'hd84;
    assign memory[6065] = 12'hd84;
    assign memory[6066] = 12'hd84;
    assign memory[6067] = 12'hd84;
    assign memory[6068] = 12'hd84;
    assign memory[6069] = 12'hd84;
    assign memory[6070] = 12'hd84;
    assign memory[6071] = 12'hd84;
    assign memory[6072] = 12'hd84;
    assign memory[6073] = 12'hd84;
    assign memory[6074] = 12'hd84;
    assign memory[6075] = 12'hd84;
    assign memory[6076] = 12'hd84;
    assign memory[6077] = 12'hd84;
    assign memory[6078] = 12'hd84;
    assign memory[6079] = 12'hc94;
    assign memory[6080] = 12'hd84;
    assign memory[6081] = 12'hd84;
    assign memory[6082] = 12'hd84;
    assign memory[6083] = 12'hd84;
    assign memory[6084] = 12'hd84;
    assign memory[6085] = 12'hd84;
    assign memory[6086] = 12'hd84;
    assign memory[6087] = 12'hd84;
    assign memory[6088] = 12'hd84;
    assign memory[6089] = 12'hc94;
    assign memory[6090] = 12'hd84;
    assign memory[6091] = 12'hd84;
    assign memory[6092] = 12'hd84;
    assign memory[6093] = 12'hc94;
    assign memory[6094] = 12'hd74;
    assign memory[6095] = 12'hc94;
    assign memory[6096] = 12'hd84;
    assign memory[6097] = 12'hd84;
    assign memory[6098] = 12'hd84;
    assign memory[6099] = 12'hd74;
    assign memory[6100] = 12'hd84;
    assign memory[6101] = 12'hd84;
    assign memory[6102] = 12'hd84;
    assign memory[6103] = 12'hd84;
    assign memory[6104] = 12'hc94;
    assign memory[6105] = 12'hd85;
    assign memory[6106] = 12'hd84;
    assign memory[6107] = 12'hd74;
    assign memory[6108] = 12'hd84;
    assign memory[6109] = 12'hd84;
    assign memory[6110] = 12'hd84;
    assign memory[6111] = 12'hd84;
    assign memory[6112] = 12'hd84;
    assign memory[6113] = 12'hd84;
    assign memory[6114] = 12'hd84;
    assign memory[6115] = 12'hd84;
    assign memory[6116] = 12'hd84;
    assign memory[6117] = 12'hd84;
    assign memory[6118] = 12'hd84;
    assign memory[6119] = 12'hd84;
    assign memory[6120] = 12'hd84;
    assign memory[6121] = 12'hd84;
    assign memory[6122] = 12'hd84;
    assign memory[6123] = 12'hd84;
    assign memory[6124] = 12'hd74;
    assign memory[6125] = 12'hd84;
    assign memory[6126] = 12'hc94;
    assign memory[6127] = 12'hd84;
    assign memory[6128] = 12'hd84;
    assign memory[6129] = 12'hd84;
    assign memory[6130] = 12'hd84;
    assign memory[6131] = 12'hd84;
    assign memory[6132] = 12'hd84;
    assign memory[6133] = 12'hd84;
    assign memory[6134] = 12'hd84;
    assign memory[6135] = 12'hd84;
    assign memory[6136] = 12'hd84;
    assign memory[6137] = 12'hd84;
    assign memory[6138] = 12'hd85;
    assign memory[6139] = 12'hd84;
    assign memory[6140] = 12'hd84;
    assign memory[6141] = 12'hd84;
    assign memory[6142] = 12'hd84;
    assign memory[6143] = 12'hd84;
    assign memory[6144] = 12'h600;
    assign memory[6145] = 12'h801;
    assign memory[6146] = 12'h901;
    assign memory[6147] = 12'h901;
    assign memory[6148] = 12'h901;
    assign memory[6149] = 12'h901;
    assign memory[6150] = 12'h901;
    assign memory[6151] = 12'h901;
    assign memory[6152] = 12'h901;
    assign memory[6153] = 12'h901;
    assign memory[6154] = 12'h901;
    assign memory[6155] = 12'h901;
    assign memory[6156] = 12'h901;
    assign memory[6157] = 12'h901;
    assign memory[6158] = 12'h901;
    assign memory[6159] = 12'h901;
    assign memory[6160] = 12'h901;
    assign memory[6161] = 12'h901;
    assign memory[6162] = 12'h901;
    assign memory[6163] = 12'h901;
    assign memory[6164] = 12'h901;
    assign memory[6165] = 12'h901;
    assign memory[6166] = 12'h901;
    assign memory[6167] = 12'h901;
    assign memory[6168] = 12'h901;
    assign memory[6169] = 12'h901;
    assign memory[6170] = 12'h901;
    assign memory[6171] = 12'h901;
    assign memory[6172] = 12'h901;
    assign memory[6173] = 12'h901;
    assign memory[6174] = 12'h801;
    assign memory[6175] = 12'h600;
    assign memory[6176] = 12'h801;
    assign memory[6177] = 12'h600;
    assign memory[6178] = 12'h801;
    assign memory[6179] = 12'h901;
    assign memory[6180] = 12'h901;
    assign memory[6181] = 12'h901;
    assign memory[6182] = 12'h901;
    assign memory[6183] = 12'h901;
    assign memory[6184] = 12'h901;
    assign memory[6185] = 12'h901;
    assign memory[6186] = 12'h901;
    assign memory[6187] = 12'h901;
    assign memory[6188] = 12'h901;
    assign memory[6189] = 12'h901;
    assign memory[6190] = 12'h901;
    assign memory[6191] = 12'h901;
    assign memory[6192] = 12'h901;
    assign memory[6193] = 12'h901;
    assign memory[6194] = 12'h901;
    assign memory[6195] = 12'h901;
    assign memory[6196] = 12'h901;
    assign memory[6197] = 12'h901;
    assign memory[6198] = 12'h901;
    assign memory[6199] = 12'h901;
    assign memory[6200] = 12'h901;
    assign memory[6201] = 12'h901;
    assign memory[6202] = 12'h901;
    assign memory[6203] = 12'h901;
    assign memory[6204] = 12'h901;
    assign memory[6205] = 12'h801;
    assign memory[6206] = 12'h600;
    assign memory[6207] = 12'h801;
    assign memory[6208] = 12'h901;
    assign memory[6209] = 12'h801;
    assign memory[6210] = 12'h600;
    assign memory[6211] = 12'h801;
    assign memory[6212] = 12'h901;
    assign memory[6213] = 12'h901;
    assign memory[6214] = 12'h901;
    assign memory[6215] = 12'h901;
    assign memory[6216] = 12'h901;
    assign memory[6217] = 12'h901;
    assign memory[6218] = 12'h901;
    assign memory[6219] = 12'h901;
    assign memory[6220] = 12'h901;
    assign memory[6221] = 12'h901;
    assign memory[6222] = 12'h901;
    assign memory[6223] = 12'h901;
    assign memory[6224] = 12'h901;
    assign memory[6225] = 12'h901;
    assign memory[6226] = 12'h901;
    assign memory[6227] = 12'h901;
    assign memory[6228] = 12'h901;
    assign memory[6229] = 12'h901;
    assign memory[6230] = 12'h901;
    assign memory[6231] = 12'h901;
    assign memory[6232] = 12'h901;
    assign memory[6233] = 12'h901;
    assign memory[6234] = 12'h901;
    assign memory[6235] = 12'h901;
    assign memory[6236] = 12'h801;
    assign memory[6237] = 12'h600;
    assign memory[6238] = 12'h801;
    assign memory[6239] = 12'h901;
    assign memory[6240] = 12'h901;
    assign memory[6241] = 12'h901;
    assign memory[6242] = 12'h801;
    assign memory[6243] = 12'h600;
    assign memory[6244] = 12'h801;
    assign memory[6245] = 12'h901;
    assign memory[6246] = 12'h901;
    assign memory[6247] = 12'h901;
    assign memory[6248] = 12'h901;
    assign memory[6249] = 12'h901;
    assign memory[6250] = 12'h901;
    assign memory[6251] = 12'h901;
    assign memory[6252] = 12'h901;
    assign memory[6253] = 12'h901;
    assign memory[6254] = 12'h901;
    assign memory[6255] = 12'h901;
    assign memory[6256] = 12'h901;
    assign memory[6257] = 12'h901;
    assign memory[6258] = 12'h901;
    assign memory[6259] = 12'h901;
    assign memory[6260] = 12'h901;
    assign memory[6261] = 12'h901;
    assign memory[6262] = 12'h901;
    assign memory[6263] = 12'h901;
    assign memory[6264] = 12'h901;
    assign memory[6265] = 12'h901;
    assign memory[6266] = 12'h901;
    assign memory[6267] = 12'h801;
    assign memory[6268] = 12'h600;
    assign memory[6269] = 12'h801;
    assign memory[6270] = 12'h901;
    assign memory[6271] = 12'h901;
    assign memory[6272] = 12'h901;
    assign memory[6273] = 12'h901;
    assign memory[6274] = 12'h901;
    assign memory[6275] = 12'h801;
    assign memory[6276] = 12'h600;
    assign memory[6277] = 12'h801;
    assign memory[6278] = 12'h901;
    assign memory[6279] = 12'h901;
    assign memory[6280] = 12'h901;
    assign memory[6281] = 12'h901;
    assign memory[6282] = 12'h901;
    assign memory[6283] = 12'h901;
    assign memory[6284] = 12'h901;
    assign memory[6285] = 12'h901;
    assign memory[6286] = 12'h901;
    assign memory[6287] = 12'h901;
    assign memory[6288] = 12'h901;
    assign memory[6289] = 12'h901;
    assign memory[6290] = 12'h901;
    assign memory[6291] = 12'h901;
    assign memory[6292] = 12'h901;
    assign memory[6293] = 12'h901;
    assign memory[6294] = 12'h901;
    assign memory[6295] = 12'h901;
    assign memory[6296] = 12'h901;
    assign memory[6297] = 12'h901;
    assign memory[6298] = 12'h801;
    assign memory[6299] = 12'h600;
    assign memory[6300] = 12'h801;
    assign memory[6301] = 12'h901;
    assign memory[6302] = 12'h901;
    assign memory[6303] = 12'h901;
    assign memory[6304] = 12'h901;
    assign memory[6305] = 12'h901;
    assign memory[6306] = 12'h901;
    assign memory[6307] = 12'h901;
    assign memory[6308] = 12'hff0;
    assign memory[6309] = 12'h600;
    assign memory[6310] = 12'h801;
    assign memory[6311] = 12'h901;
    assign memory[6312] = 12'h901;
    assign memory[6313] = 12'h901;
    assign memory[6314] = 12'h901;
    assign memory[6315] = 12'h901;
    assign memory[6316] = 12'h901;
    assign memory[6317] = 12'h901;
    assign memory[6318] = 12'h901;
    assign memory[6319] = 12'h901;
    assign memory[6320] = 12'h901;
    assign memory[6321] = 12'h901;
    assign memory[6322] = 12'h901;
    assign memory[6323] = 12'h901;
    assign memory[6324] = 12'h901;
    assign memory[6325] = 12'h901;
    assign memory[6326] = 12'h901;
    assign memory[6327] = 12'h901;
    assign memory[6328] = 12'h901;
    assign memory[6329] = 12'h801;
    assign memory[6330] = 12'h600;
    assign memory[6331] = 12'h801;
    assign memory[6332] = 12'h901;
    assign memory[6333] = 12'h901;
    assign memory[6334] = 12'h901;
    assign memory[6335] = 12'h901;
    assign memory[6336] = 12'h901;
    assign memory[6337] = 12'hccc;
    assign memory[6338] = 12'h901;
    assign memory[6339] = 12'hff0;
    assign memory[6340] = 12'hff0;
    assign memory[6341] = 12'h901;
    assign memory[6342] = 12'hccc;
    assign memory[6343] = 12'h801;
    assign memory[6344] = 12'h901;
    assign memory[6345] = 12'h901;
    assign memory[6346] = 12'h901;
    assign memory[6347] = 12'h901;
    assign memory[6348] = 12'h901;
    assign memory[6349] = 12'h901;
    assign memory[6350] = 12'h901;
    assign memory[6351] = 12'h901;
    assign memory[6352] = 12'h901;
    assign memory[6353] = 12'h901;
    assign memory[6354] = 12'h901;
    assign memory[6355] = 12'h901;
    assign memory[6356] = 12'h901;
    assign memory[6357] = 12'h901;
    assign memory[6358] = 12'h901;
    assign memory[6359] = 12'h901;
    assign memory[6360] = 12'h801;
    assign memory[6361] = 12'h600;
    assign memory[6362] = 12'h801;
    assign memory[6363] = 12'h901;
    assign memory[6364] = 12'h901;
    assign memory[6365] = 12'h901;
    assign memory[6366] = 12'h901;
    assign memory[6367] = 12'h901;
    assign memory[6368] = 12'h901;
    assign memory[6369] = 12'hccc;
    assign memory[6370] = 12'h901;
    assign memory[6371] = 12'hff0;
    assign memory[6372] = 12'hff0;
    assign memory[6373] = 12'h901;
    assign memory[6374] = 12'hccc;
    assign memory[6375] = 12'h600;
    assign memory[6376] = 12'h801;
    assign memory[6377] = 12'h901;
    assign memory[6378] = 12'h901;
    assign memory[6379] = 12'h901;
    assign memory[6380] = 12'h901;
    assign memory[6381] = 12'h901;
    assign memory[6382] = 12'h901;
    assign memory[6383] = 12'h901;
    assign memory[6384] = 12'h901;
    assign memory[6385] = 12'h901;
    assign memory[6386] = 12'h901;
    assign memory[6387] = 12'h901;
    assign memory[6388] = 12'h901;
    assign memory[6389] = 12'h901;
    assign memory[6390] = 12'h901;
    assign memory[6391] = 12'h801;
    assign memory[6392] = 12'h600;
    assign memory[6393] = 12'h801;
    assign memory[6394] = 12'h901;
    assign memory[6395] = 12'h901;
    assign memory[6396] = 12'h901;
    assign memory[6397] = 12'h901;
    assign memory[6398] = 12'h901;
    assign memory[6399] = 12'h901;
    assign memory[6400] = 12'h901;
    assign memory[6401] = 12'hccc;
    assign memory[6402] = 12'hffd;
    assign memory[6403] = 12'hffd;
    assign memory[6404] = 12'hffd;
    assign memory[6405] = 12'hffd;
    assign memory[6406] = 12'hccc;
    assign memory[6407] = 12'h801;
    assign memory[6408] = 12'h600;
    assign memory[6409] = 12'h801;
    assign memory[6410] = 12'h901;
    assign memory[6411] = 12'h901;
    assign memory[6412] = 12'h901;
    assign memory[6413] = 12'h901;
    assign memory[6414] = 12'h901;
    assign memory[6415] = 12'h901;
    assign memory[6416] = 12'h901;
    assign memory[6417] = 12'h901;
    assign memory[6418] = 12'h901;
    assign memory[6419] = 12'h901;
    assign memory[6420] = 12'h901;
    assign memory[6421] = 12'h901;
    assign memory[6422] = 12'h801;
    assign memory[6423] = 12'h600;
    assign memory[6424] = 12'h801;
    assign memory[6425] = 12'h901;
    assign memory[6426] = 12'h901;
    assign memory[6427] = 12'h901;
    assign memory[6428] = 12'h901;
    assign memory[6429] = 12'h901;
    assign memory[6430] = 12'h901;
    assign memory[6431] = 12'h901;
    assign memory[6432] = 12'h901;
    assign memory[6433] = 12'hccc;
    assign memory[6434] = 12'hffd;
    assign memory[6435] = 12'hffd;
    assign memory[6436] = 12'hffd;
    assign memory[6437] = 12'hffd;
    assign memory[6438] = 12'hccc;
    assign memory[6439] = 12'h901;
    assign memory[6440] = 12'h801;
    assign memory[6441] = 12'h600;
    assign memory[6442] = 12'h801;
    assign memory[6443] = 12'h901;
    assign memory[6444] = 12'h901;
    assign memory[6445] = 12'h901;
    assign memory[6446] = 12'h901;
    assign memory[6447] = 12'h901;
    assign memory[6448] = 12'h901;
    assign memory[6449] = 12'h901;
    assign memory[6450] = 12'h901;
    assign memory[6451] = 12'h901;
    assign memory[6452] = 12'h901;
    assign memory[6453] = 12'h801;
    assign memory[6454] = 12'h600;
    assign memory[6455] = 12'h801;
    assign memory[6456] = 12'h901;
    assign memory[6457] = 12'h901;
    assign memory[6458] = 12'h901;
    assign memory[6459] = 12'h901;
    assign memory[6460] = 12'h901;
    assign memory[6461] = 12'h901;
    assign memory[6462] = 12'h901;
    assign memory[6463] = 12'h901;
    assign memory[6464] = 12'h901;
    assign memory[6465] = 12'hccc;
    assign memory[6466] = 12'hffd;
    assign memory[6467] = 12'hffd;
    assign memory[6468] = 12'hffd;
    assign memory[6469] = 12'hffd;
    assign memory[6470] = 12'hccc;
    assign memory[6471] = 12'h901;
    assign memory[6472] = 12'h901;
    assign memory[6473] = 12'h801;
    assign memory[6474] = 12'h600;
    assign memory[6475] = 12'h801;
    assign memory[6476] = 12'h901;
    assign memory[6477] = 12'h901;
    assign memory[6478] = 12'h901;
    assign memory[6479] = 12'h901;
    assign memory[6480] = 12'h901;
    assign memory[6481] = 12'h901;
    assign memory[6482] = 12'h901;
    assign memory[6483] = 12'h901;
    assign memory[6484] = 12'h801;
    assign memory[6485] = 12'h600;
    assign memory[6486] = 12'h801;
    assign memory[6487] = 12'h901;
    assign memory[6488] = 12'h901;
    assign memory[6489] = 12'h901;
    assign memory[6490] = 12'h901;
    assign memory[6491] = 12'h901;
    assign memory[6492] = 12'h901;
    assign memory[6493] = 12'h901;
    assign memory[6494] = 12'h901;
    assign memory[6495] = 12'h901;
    assign memory[6496] = 12'h901;
    assign memory[6497] = 12'hccc;
    assign memory[6498] = 12'hffd;
    assign memory[6499] = 12'hffd;
    assign memory[6500] = 12'hffd;
    assign memory[6501] = 12'hffd;
    assign memory[6502] = 12'hccc;
    assign memory[6503] = 12'h901;
    assign memory[6504] = 12'h901;
    assign memory[6505] = 12'h901;
    assign memory[6506] = 12'h801;
    assign memory[6507] = 12'h600;
    assign memory[6508] = 12'h801;
    assign memory[6509] = 12'h901;
    assign memory[6510] = 12'h901;
    assign memory[6511] = 12'h901;
    assign memory[6512] = 12'h901;
    assign memory[6513] = 12'h901;
    assign memory[6514] = 12'h901;
    assign memory[6515] = 12'h801;
    assign memory[6516] = 12'h600;
    assign memory[6517] = 12'h801;
    assign memory[6518] = 12'h901;
    assign memory[6519] = 12'h901;
    assign memory[6520] = 12'h901;
    assign memory[6521] = 12'h901;
    assign memory[6522] = 12'h901;
    assign memory[6523] = 12'h901;
    assign memory[6524] = 12'h901;
    assign memory[6525] = 12'h901;
    assign memory[6526] = 12'h901;
    assign memory[6527] = 12'h901;
    assign memory[6528] = 12'h901;
    assign memory[6529] = 12'hccc;
    assign memory[6530] = 12'hccc;
    assign memory[6531] = 12'hccc;
    assign memory[6532] = 12'hccc;
    assign memory[6533] = 12'hccc;
    assign memory[6534] = 12'hccc;
    assign memory[6535] = 12'h901;
    assign memory[6536] = 12'h901;
    assign memory[6537] = 12'h901;
    assign memory[6538] = 12'h901;
    assign memory[6539] = 12'h801;
    assign memory[6540] = 12'h600;
    assign memory[6541] = 12'h801;
    assign memory[6542] = 12'h901;
    assign memory[6543] = 12'h901;
    assign memory[6544] = 12'h901;
    assign memory[6545] = 12'h901;
    assign memory[6546] = 12'h801;
    assign memory[6547] = 12'h600;
    assign memory[6548] = 12'h801;
    assign memory[6549] = 12'h901;
    assign memory[6550] = 12'h901;
    assign memory[6551] = 12'h901;
    assign memory[6552] = 12'h901;
    assign memory[6553] = 12'h901;
    assign memory[6554] = 12'h901;
    assign memory[6555] = 12'h901;
    assign memory[6556] = 12'h901;
    assign memory[6557] = 12'h901;
    assign memory[6558] = 12'h901;
    assign memory[6559] = 12'h901;
    assign memory[6560] = 12'h901;
    assign memory[6561] = 12'h901;
    assign memory[6562] = 12'h901;
    assign memory[6563] = 12'h901;
    assign memory[6564] = 12'h901;
    assign memory[6565] = 12'h901;
    assign memory[6566] = 12'h901;
    assign memory[6567] = 12'h901;
    assign memory[6568] = 12'h901;
    assign memory[6569] = 12'h901;
    assign memory[6570] = 12'h901;
    assign memory[6571] = 12'h901;
    assign memory[6572] = 12'h801;
    assign memory[6573] = 12'h600;
    assign memory[6574] = 12'h801;
    assign memory[6575] = 12'h901;
    assign memory[6576] = 12'h901;
    assign memory[6577] = 12'h801;
    assign memory[6578] = 12'h600;
    assign memory[6579] = 12'h801;
    assign memory[6580] = 12'h901;
    assign memory[6581] = 12'h901;
    assign memory[6582] = 12'h901;
    assign memory[6583] = 12'h901;
    assign memory[6584] = 12'h901;
    assign memory[6585] = 12'h901;
    assign memory[6586] = 12'h901;
    assign memory[6587] = 12'h901;
    assign memory[6588] = 12'h901;
    assign memory[6589] = 12'h901;
    assign memory[6590] = 12'h901;
    assign memory[6591] = 12'h901;
    assign memory[6592] = 12'h901;
    assign memory[6593] = 12'h901;
    assign memory[6594] = 12'h901;
    assign memory[6595] = 12'h901;
    assign memory[6596] = 12'h901;
    assign memory[6597] = 12'h901;
    assign memory[6598] = 12'h901;
    assign memory[6599] = 12'h901;
    assign memory[6600] = 12'h901;
    assign memory[6601] = 12'h901;
    assign memory[6602] = 12'h901;
    assign memory[6603] = 12'h901;
    assign memory[6604] = 12'h901;
    assign memory[6605] = 12'h801;
    assign memory[6606] = 12'h600;
    assign memory[6607] = 12'h801;
    assign memory[6608] = 12'h801;
    assign memory[6609] = 12'h600;
    assign memory[6610] = 12'h801;
    assign memory[6611] = 12'h901;
    assign memory[6612] = 12'h901;
    assign memory[6613] = 12'h901;
    assign memory[6614] = 12'h901;
    assign memory[6615] = 12'h901;
    assign memory[6616] = 12'h901;
    assign memory[6617] = 12'h901;
    assign memory[6618] = 12'h901;
    assign memory[6619] = 12'h901;
    assign memory[6620] = 12'h901;
    assign memory[6621] = 12'h901;
    assign memory[6622] = 12'h901;
    assign memory[6623] = 12'h901;
    assign memory[6624] = 12'h901;
    assign memory[6625] = 12'h901;
    assign memory[6626] = 12'h901;
    assign memory[6627] = 12'h901;
    assign memory[6628] = 12'h901;
    assign memory[6629] = 12'h901;
    assign memory[6630] = 12'h901;
    assign memory[6631] = 12'h901;
    assign memory[6632] = 12'h901;
    assign memory[6633] = 12'h901;
    assign memory[6634] = 12'h901;
    assign memory[6635] = 12'h901;
    assign memory[6636] = 12'h901;
    assign memory[6637] = 12'h901;
    assign memory[6638] = 12'h801;
    assign memory[6639] = 12'h600;
    assign memory[6640] = 12'h600;
    assign memory[6641] = 12'h801;
    assign memory[6642] = 12'h901;
    assign memory[6643] = 12'h901;
    assign memory[6644] = 12'h901;
    assign memory[6645] = 12'h901;
    assign memory[6646] = 12'h901;
    assign memory[6647] = 12'h901;
    assign memory[6648] = 12'h901;
    assign memory[6649] = 12'h901;
    assign memory[6650] = 12'h901;
    assign memory[6651] = 12'h901;
    assign memory[6652] = 12'h901;
    assign memory[6653] = 12'h901;
    assign memory[6654] = 12'h901;
    assign memory[6655] = 12'h901;
    assign memory[6656] = 12'h901;
    assign memory[6657] = 12'h901;
    assign memory[6658] = 12'h901;
    assign memory[6659] = 12'h901;
    assign memory[6660] = 12'h901;
    assign memory[6661] = 12'h901;
    assign memory[6662] = 12'h901;
    assign memory[6663] = 12'h901;
    assign memory[6664] = 12'h901;
    assign memory[6665] = 12'h901;
    assign memory[6666] = 12'h901;
    assign memory[6667] = 12'h901;
    assign memory[6668] = 12'h901;
    assign memory[6669] = 12'h901;
    assign memory[6670] = 12'h801;
    assign memory[6671] = 12'h600;
    assign memory[6672] = 12'h600;
    assign memory[6673] = 12'h801;
    assign memory[6674] = 12'h901;
    assign memory[6675] = 12'h901;
    assign memory[6676] = 12'h901;
    assign memory[6677] = 12'h901;
    assign memory[6678] = 12'h901;
    assign memory[6679] = 12'h901;
    assign memory[6680] = 12'h901;
    assign memory[6681] = 12'h901;
    assign memory[6682] = 12'h901;
    assign memory[6683] = 12'h901;
    assign memory[6684] = 12'h901;
    assign memory[6685] = 12'h901;
    assign memory[6686] = 12'h901;
    assign memory[6687] = 12'h901;
    assign memory[6688] = 12'h901;
    assign memory[6689] = 12'h901;
    assign memory[6690] = 12'h901;
    assign memory[6691] = 12'h901;
    assign memory[6692] = 12'h901;
    assign memory[6693] = 12'h901;
    assign memory[6694] = 12'h901;
    assign memory[6695] = 12'h901;
    assign memory[6696] = 12'h901;
    assign memory[6697] = 12'h901;
    assign memory[6698] = 12'h901;
    assign memory[6699] = 12'h901;
    assign memory[6700] = 12'h901;
    assign memory[6701] = 12'h801;
    assign memory[6702] = 12'h600;
    assign memory[6703] = 12'h801;
    assign memory[6704] = 12'h801;
    assign memory[6705] = 12'h600;
    assign memory[6706] = 12'h801;
    assign memory[6707] = 12'h901;
    assign memory[6708] = 12'h901;
    assign memory[6709] = 12'h901;
    assign memory[6710] = 12'h901;
    assign memory[6711] = 12'h901;
    assign memory[6712] = 12'h901;
    assign memory[6713] = 12'h901;
    assign memory[6714] = 12'h901;
    assign memory[6715] = 12'h901;
    assign memory[6716] = 12'h901;
    assign memory[6717] = 12'h901;
    assign memory[6718] = 12'h901;
    assign memory[6719] = 12'h901;
    assign memory[6720] = 12'h901;
    assign memory[6721] = 12'h901;
    assign memory[6722] = 12'h901;
    assign memory[6723] = 12'h901;
    assign memory[6724] = 12'h901;
    assign memory[6725] = 12'h901;
    assign memory[6726] = 12'h901;
    assign memory[6727] = 12'h901;
    assign memory[6728] = 12'h901;
    assign memory[6729] = 12'h901;
    assign memory[6730] = 12'h901;
    assign memory[6731] = 12'h901;
    assign memory[6732] = 12'h801;
    assign memory[6733] = 12'h600;
    assign memory[6734] = 12'h801;
    assign memory[6735] = 12'h901;
    assign memory[6736] = 12'h901;
    assign memory[6737] = 12'h801;
    assign memory[6738] = 12'h600;
    assign memory[6739] = 12'h801;
    assign memory[6740] = 12'h901;
    assign memory[6741] = 12'h901;
    assign memory[6742] = 12'h901;
    assign memory[6743] = 12'h901;
    assign memory[6744] = 12'h901;
    assign memory[6745] = 12'h901;
    assign memory[6746] = 12'h901;
    assign memory[6747] = 12'h901;
    assign memory[6748] = 12'h901;
    assign memory[6749] = 12'h901;
    assign memory[6750] = 12'h901;
    assign memory[6751] = 12'h901;
    assign memory[6752] = 12'h901;
    assign memory[6753] = 12'h901;
    assign memory[6754] = 12'h901;
    assign memory[6755] = 12'h901;
    assign memory[6756] = 12'h901;
    assign memory[6757] = 12'h901;
    assign memory[6758] = 12'h901;
    assign memory[6759] = 12'h901;
    assign memory[6760] = 12'h901;
    assign memory[6761] = 12'h901;
    assign memory[6762] = 12'h901;
    assign memory[6763] = 12'h801;
    assign memory[6764] = 12'h600;
    assign memory[6765] = 12'h801;
    assign memory[6766] = 12'h901;
    assign memory[6767] = 12'h901;
    assign memory[6768] = 12'h901;
    assign memory[6769] = 12'h901;
    assign memory[6770] = 12'h801;
    assign memory[6771] = 12'h600;
    assign memory[6772] = 12'h801;
    assign memory[6773] = 12'h901;
    assign memory[6774] = 12'h901;
    assign memory[6775] = 12'h901;
    assign memory[6776] = 12'h901;
    assign memory[6777] = 12'h901;
    assign memory[6778] = 12'h901;
    assign memory[6779] = 12'h901;
    assign memory[6780] = 12'h901;
    assign memory[6781] = 12'h901;
    assign memory[6782] = 12'h901;
    assign memory[6783] = 12'h901;
    assign memory[6784] = 12'h901;
    assign memory[6785] = 12'h901;
    assign memory[6786] = 12'h901;
    assign memory[6787] = 12'h901;
    assign memory[6788] = 12'h901;
    assign memory[6789] = 12'h901;
    assign memory[6790] = 12'h901;
    assign memory[6791] = 12'h901;
    assign memory[6792] = 12'h901;
    assign memory[6793] = 12'h901;
    assign memory[6794] = 12'h801;
    assign memory[6795] = 12'h600;
    assign memory[6796] = 12'h801;
    assign memory[6797] = 12'h901;
    assign memory[6798] = 12'h901;
    assign memory[6799] = 12'h901;
    assign memory[6800] = 12'h901;
    assign memory[6801] = 12'h901;
    assign memory[6802] = 12'h901;
    assign memory[6803] = 12'h801;
    assign memory[6804] = 12'h600;
    assign memory[6805] = 12'h801;
    assign memory[6806] = 12'h901;
    assign memory[6807] = 12'h901;
    assign memory[6808] = 12'h901;
    assign memory[6809] = 12'h901;
    assign memory[6810] = 12'h901;
    assign memory[6811] = 12'h901;
    assign memory[6812] = 12'h901;
    assign memory[6813] = 12'h901;
    assign memory[6814] = 12'h901;
    assign memory[6815] = 12'h901;
    assign memory[6816] = 12'h901;
    assign memory[6817] = 12'h901;
    assign memory[6818] = 12'h901;
    assign memory[6819] = 12'h901;
    assign memory[6820] = 12'h901;
    assign memory[6821] = 12'h901;
    assign memory[6822] = 12'h901;
    assign memory[6823] = 12'h901;
    assign memory[6824] = 12'h901;
    assign memory[6825] = 12'h801;
    assign memory[6826] = 12'h600;
    assign memory[6827] = 12'h801;
    assign memory[6828] = 12'h901;
    assign memory[6829] = 12'h901;
    assign memory[6830] = 12'h901;
    assign memory[6831] = 12'h901;
    assign memory[6832] = 12'h901;
    assign memory[6833] = 12'h901;
    assign memory[6834] = 12'h901;
    assign memory[6835] = 12'h901;
    assign memory[6836] = 12'h801;
    assign memory[6837] = 12'h600;
    assign memory[6838] = 12'h901;
    assign memory[6839] = 12'h901;
    assign memory[6840] = 12'h901;
    assign memory[6841] = 12'h901;
    assign memory[6842] = 12'h901;
    assign memory[6843] = 12'h901;
    assign memory[6844] = 12'h901;
    assign memory[6845] = 12'h901;
    assign memory[6846] = 12'h901;
    assign memory[6847] = 12'h901;
    assign memory[6848] = 12'h901;
    assign memory[6849] = 12'h901;
    assign memory[6850] = 12'h901;
    assign memory[6851] = 12'h901;
    assign memory[6852] = 12'h901;
    assign memory[6853] = 12'h901;
    assign memory[6854] = 12'h901;
    assign memory[6855] = 12'h901;
    assign memory[6856] = 12'h801;
    assign memory[6857] = 12'h600;
    assign memory[6858] = 12'h801;
    assign memory[6859] = 12'h901;
    assign memory[6860] = 12'h901;
    assign memory[6861] = 12'h901;
    assign memory[6862] = 12'h901;
    assign memory[6863] = 12'h901;
    assign memory[6864] = 12'h901;
    assign memory[6865] = 12'h901;
    assign memory[6866] = 12'h901;
    assign memory[6867] = 12'h901;
    assign memory[6868] = 12'h901;
    assign memory[6869] = 12'h801;
    assign memory[6870] = 12'h600;
    assign memory[6871] = 12'h801;
    assign memory[6872] = 12'h901;
    assign memory[6873] = 12'h901;
    assign memory[6874] = 12'h901;
    assign memory[6875] = 12'h901;
    assign memory[6876] = 12'h901;
    assign memory[6877] = 12'h901;
    assign memory[6878] = 12'h901;
    assign memory[6879] = 12'h901;
    assign memory[6880] = 12'h901;
    assign memory[6881] = 12'h901;
    assign memory[6882] = 12'h901;
    assign memory[6883] = 12'h901;
    assign memory[6884] = 12'h901;
    assign memory[6885] = 12'h901;
    assign memory[6886] = 12'h901;
    assign memory[6887] = 12'h801;
    assign memory[6888] = 12'h600;
    assign memory[6889] = 12'h801;
    assign memory[6890] = 12'h901;
    assign memory[6891] = 12'h901;
    assign memory[6892] = 12'h901;
    assign memory[6893] = 12'h901;
    assign memory[6894] = 12'h901;
    assign memory[6895] = 12'h901;
    assign memory[6896] = 12'h901;
    assign memory[6897] = 12'h901;
    assign memory[6898] = 12'h901;
    assign memory[6899] = 12'h901;
    assign memory[6900] = 12'h901;
    assign memory[6901] = 12'h901;
    assign memory[6902] = 12'h801;
    assign memory[6903] = 12'h600;
    assign memory[6904] = 12'h801;
    assign memory[6905] = 12'h901;
    assign memory[6906] = 12'h901;
    assign memory[6907] = 12'h901;
    assign memory[6908] = 12'h901;
    assign memory[6909] = 12'h901;
    assign memory[6910] = 12'h901;
    assign memory[6911] = 12'h901;
    assign memory[6912] = 12'h901;
    assign memory[6913] = 12'h901;
    assign memory[6914] = 12'h901;
    assign memory[6915] = 12'h901;
    assign memory[6916] = 12'h901;
    assign memory[6917] = 12'h901;
    assign memory[6918] = 12'h801;
    assign memory[6919] = 12'h600;
    assign memory[6920] = 12'h801;
    assign memory[6921] = 12'h901;
    assign memory[6922] = 12'h901;
    assign memory[6923] = 12'h901;
    assign memory[6924] = 12'h901;
    assign memory[6925] = 12'h901;
    assign memory[6926] = 12'h901;
    assign memory[6927] = 12'h901;
    assign memory[6928] = 12'h901;
    assign memory[6929] = 12'h901;
    assign memory[6930] = 12'h901;
    assign memory[6931] = 12'h901;
    assign memory[6932] = 12'h901;
    assign memory[6933] = 12'h901;
    assign memory[6934] = 12'h901;
    assign memory[6935] = 12'h801;
    assign memory[6936] = 12'h600;
    assign memory[6937] = 12'hff0;
    assign memory[6938] = 12'h901;
    assign memory[6939] = 12'h901;
    assign memory[6940] = 12'h901;
    assign memory[6941] = 12'h901;
    assign memory[6942] = 12'h901;
    assign memory[6943] = 12'h901;
    assign memory[6944] = 12'h901;
    assign memory[6945] = 12'h901;
    assign memory[6946] = 12'h901;
    assign memory[6947] = 12'h901;
    assign memory[6948] = 12'h901;
    assign memory[6949] = 12'h801;
    assign memory[6950] = 12'h600;
    assign memory[6951] = 12'h801;
    assign memory[6952] = 12'h901;
    assign memory[6953] = 12'h901;
    assign memory[6954] = 12'h901;
    assign memory[6955] = 12'h901;
    assign memory[6956] = 12'h901;
    assign memory[6957] = 12'h901;
    assign memory[6958] = 12'h901;
    assign memory[6959] = 12'h901;
    assign memory[6960] = 12'h901;
    assign memory[6961] = 12'h901;
    assign memory[6962] = 12'h901;
    assign memory[6963] = 12'h901;
    assign memory[6964] = 12'h901;
    assign memory[6965] = 12'h901;
    assign memory[6966] = 12'hccc;
    assign memory[6967] = 12'h901;
    assign memory[6968] = 12'hff0;
    assign memory[6969] = 12'hff0;
    assign memory[6970] = 12'h901;
    assign memory[6971] = 12'hccc;
    assign memory[6972] = 12'h901;
    assign memory[6973] = 12'h901;
    assign memory[6974] = 12'h901;
    assign memory[6975] = 12'h901;
    assign memory[6976] = 12'h901;
    assign memory[6977] = 12'h901;
    assign memory[6978] = 12'h901;
    assign memory[6979] = 12'h901;
    assign memory[6980] = 12'h801;
    assign memory[6981] = 12'h600;
    assign memory[6982] = 12'h801;
    assign memory[6983] = 12'h901;
    assign memory[6984] = 12'h901;
    assign memory[6985] = 12'h901;
    assign memory[6986] = 12'h901;
    assign memory[6987] = 12'h901;
    assign memory[6988] = 12'h901;
    assign memory[6989] = 12'h901;
    assign memory[6990] = 12'h901;
    assign memory[6991] = 12'h901;
    assign memory[6992] = 12'h901;
    assign memory[6993] = 12'h901;
    assign memory[6994] = 12'h901;
    assign memory[6995] = 12'h901;
    assign memory[6996] = 12'h901;
    assign memory[6997] = 12'h901;
    assign memory[6998] = 12'hccc;
    assign memory[6999] = 12'h901;
    assign memory[7000] = 12'hff0;
    assign memory[7001] = 12'hff0;
    assign memory[7002] = 12'h600;
    assign memory[7003] = 12'hccc;
    assign memory[7004] = 12'h901;
    assign memory[7005] = 12'h901;
    assign memory[7006] = 12'h901;
    assign memory[7007] = 12'h901;
    assign memory[7008] = 12'h901;
    assign memory[7009] = 12'h901;
    assign memory[7010] = 12'h901;
    assign memory[7011] = 12'h801;
    assign memory[7012] = 12'h600;
    assign memory[7013] = 12'h801;
    assign memory[7014] = 12'h901;
    assign memory[7015] = 12'h901;
    assign memory[7016] = 12'h901;
    assign memory[7017] = 12'h901;
    assign memory[7018] = 12'h901;
    assign memory[7019] = 12'h901;
    assign memory[7020] = 12'h901;
    assign memory[7021] = 12'h901;
    assign memory[7022] = 12'h901;
    assign memory[7023] = 12'h901;
    assign memory[7024] = 12'h901;
    assign memory[7025] = 12'h901;
    assign memory[7026] = 12'h901;
    assign memory[7027] = 12'h901;
    assign memory[7028] = 12'h901;
    assign memory[7029] = 12'h901;
    assign memory[7030] = 12'hccc;
    assign memory[7031] = 12'hffd;
    assign memory[7032] = 12'hffd;
    assign memory[7033] = 12'hffd;
    assign memory[7034] = 12'hffd;
    assign memory[7035] = 12'hccc;
    assign memory[7036] = 12'h801;
    assign memory[7037] = 12'h901;
    assign memory[7038] = 12'h901;
    assign memory[7039] = 12'h901;
    assign memory[7040] = 12'h901;
    assign memory[7041] = 12'h901;
    assign memory[7042] = 12'h801;
    assign memory[7043] = 12'h600;
    assign memory[7044] = 12'h801;
    assign memory[7045] = 12'h901;
    assign memory[7046] = 12'h901;
    assign memory[7047] = 12'h901;
    assign memory[7048] = 12'h901;
    assign memory[7049] = 12'h901;
    assign memory[7050] = 12'h901;
    assign memory[7051] = 12'h901;
    assign memory[7052] = 12'h901;
    assign memory[7053] = 12'h901;
    assign memory[7054] = 12'h901;
    assign memory[7055] = 12'h901;
    assign memory[7056] = 12'h901;
    assign memory[7057] = 12'h901;
    assign memory[7058] = 12'h901;
    assign memory[7059] = 12'h901;
    assign memory[7060] = 12'h901;
    assign memory[7061] = 12'h901;
    assign memory[7062] = 12'hccc;
    assign memory[7063] = 12'hffd;
    assign memory[7064] = 12'hffd;
    assign memory[7065] = 12'hffd;
    assign memory[7066] = 12'hffd;
    assign memory[7067] = 12'hccc;
    assign memory[7068] = 12'h600;
    assign memory[7069] = 12'h801;
    assign memory[7070] = 12'h901;
    assign memory[7071] = 12'h901;
    assign memory[7072] = 12'h901;
    assign memory[7073] = 12'h801;
    assign memory[7074] = 12'h600;
    assign memory[7075] = 12'h801;
    assign memory[7076] = 12'h901;
    assign memory[7077] = 12'h901;
    assign memory[7078] = 12'h901;
    assign memory[7079] = 12'h901;
    assign memory[7080] = 12'h901;
    assign memory[7081] = 12'h901;
    assign memory[7082] = 12'h901;
    assign memory[7083] = 12'h901;
    assign memory[7084] = 12'h901;
    assign memory[7085] = 12'h901;
    assign memory[7086] = 12'h901;
    assign memory[7087] = 12'h901;
    assign memory[7088] = 12'h901;
    assign memory[7089] = 12'h901;
    assign memory[7090] = 12'h901;
    assign memory[7091] = 12'h901;
    assign memory[7092] = 12'h901;
    assign memory[7093] = 12'h901;
    assign memory[7094] = 12'hccc;
    assign memory[7095] = 12'hffd;
    assign memory[7096] = 12'hffd;
    assign memory[7097] = 12'hffd;
    assign memory[7098] = 12'hffd;
    assign memory[7099] = 12'hccc;
    assign memory[7100] = 12'h801;
    assign memory[7101] = 12'h600;
    assign memory[7102] = 12'h801;
    assign memory[7103] = 12'h901;
    assign memory[7104] = 12'h801;
    assign memory[7105] = 12'h600;
    assign memory[7106] = 12'h801;
    assign memory[7107] = 12'h901;
    assign memory[7108] = 12'h901;
    assign memory[7109] = 12'h901;
    assign memory[7110] = 12'h901;
    assign memory[7111] = 12'h901;
    assign memory[7112] = 12'h901;
    assign memory[7113] = 12'h901;
    assign memory[7114] = 12'h901;
    assign memory[7115] = 12'h901;
    assign memory[7116] = 12'h901;
    assign memory[7117] = 12'h901;
    assign memory[7118] = 12'h901;
    assign memory[7119] = 12'h901;
    assign memory[7120] = 12'h901;
    assign memory[7121] = 12'h901;
    assign memory[7122] = 12'h901;
    assign memory[7123] = 12'h901;
    assign memory[7124] = 12'h901;
    assign memory[7125] = 12'h901;
    assign memory[7126] = 12'hccc;
    assign memory[7127] = 12'hffd;
    assign memory[7128] = 12'hffd;
    assign memory[7129] = 12'hffd;
    assign memory[7130] = 12'hffd;
    assign memory[7131] = 12'hccc;
    assign memory[7132] = 12'h901;
    assign memory[7133] = 12'h801;
    assign memory[7134] = 12'h600;
    assign memory[7135] = 12'h801;
    assign memory[7136] = 12'h600;
    assign memory[7137] = 12'h801;
    assign memory[7138] = 12'h901;
    assign memory[7139] = 12'h901;
    assign memory[7140] = 12'h901;
    assign memory[7141] = 12'h901;
    assign memory[7142] = 12'h901;
    assign memory[7143] = 12'h901;
    assign memory[7144] = 12'h901;
    assign memory[7145] = 12'h901;
    assign memory[7146] = 12'h901;
    assign memory[7147] = 12'h901;
    assign memory[7148] = 12'h901;
    assign memory[7149] = 12'h901;
    assign memory[7150] = 12'h901;
    assign memory[7151] = 12'h901;
    assign memory[7152] = 12'h901;
    assign memory[7153] = 12'h901;
    assign memory[7154] = 12'h901;
    assign memory[7155] = 12'h901;
    assign memory[7156] = 12'h901;
    assign memory[7157] = 12'h901;
    assign memory[7158] = 12'hccc;
    assign memory[7159] = 12'hccc;
    assign memory[7160] = 12'hccc;
    assign memory[7161] = 12'hccc;
    assign memory[7162] = 12'hccc;
    assign memory[7163] = 12'hccc;
    assign memory[7164] = 12'h901;
    assign memory[7165] = 12'h901;
    assign memory[7166] = 12'h801;
    assign memory[7167] = 12'h600;
    assign memory[7168] = 12'h654;
    assign memory[7169] = 12'h654;
    assign memory[7170] = 12'h654;
    assign memory[7171] = 12'h654;
    assign memory[7172] = 12'h654;
    assign memory[7173] = 12'h654;
    assign memory[7174] = 12'h654;
    assign memory[7175] = 12'h654;
    assign memory[7176] = 12'h654;
    assign memory[7177] = 12'h654;
    assign memory[7178] = 12'h654;
    assign memory[7179] = 12'h654;
    assign memory[7180] = 12'h654;
    assign memory[7181] = 12'h654;
    assign memory[7182] = 12'h654;
    assign memory[7183] = 12'h654;
    assign memory[7184] = 12'h654;
    assign memory[7185] = 12'h654;
    assign memory[7186] = 12'h654;
    assign memory[7187] = 12'h654;
    assign memory[7188] = 12'h654;
    assign memory[7189] = 12'h654;
    assign memory[7190] = 12'h654;
    assign memory[7191] = 12'h654;
    assign memory[7192] = 12'h654;
    assign memory[7193] = 12'h654;
    assign memory[7194] = 12'h654;
    assign memory[7195] = 12'h654;
    assign memory[7196] = 12'h654;
    assign memory[7197] = 12'h654;
    assign memory[7198] = 12'h654;
    assign memory[7199] = 12'h654;
    assign memory[7200] = 12'h654;
    assign memory[7201] = 12'h898;
    assign memory[7202] = 12'h898;
    assign memory[7203] = 12'h898;
    assign memory[7204] = 12'h898;
    assign memory[7205] = 12'h898;
    assign memory[7206] = 12'h898;
    assign memory[7207] = 12'h898;
    assign memory[7208] = 12'h898;
    assign memory[7209] = 12'h898;
    assign memory[7210] = 12'h898;
    assign memory[7211] = 12'h898;
    assign memory[7212] = 12'h898;
    assign memory[7213] = 12'h898;
    assign memory[7214] = 12'h898;
    assign memory[7215] = 12'h898;
    assign memory[7216] = 12'h898;
    assign memory[7217] = 12'h898;
    assign memory[7218] = 12'h898;
    assign memory[7219] = 12'h898;
    assign memory[7220] = 12'h898;
    assign memory[7221] = 12'h898;
    assign memory[7222] = 12'h898;
    assign memory[7223] = 12'h898;
    assign memory[7224] = 12'h898;
    assign memory[7225] = 12'h898;
    assign memory[7226] = 12'h898;
    assign memory[7227] = 12'h898;
    assign memory[7228] = 12'h898;
    assign memory[7229] = 12'h898;
    assign memory[7230] = 12'h898;
    assign memory[7231] = 12'h654;
    assign memory[7232] = 12'h654;
    assign memory[7233] = 12'h898;
    assign memory[7234] = 12'h898;
    assign memory[7235] = 12'h898;
    assign memory[7236] = 12'h898;
    assign memory[7237] = 12'h898;
    assign memory[7238] = 12'h898;
    assign memory[7239] = 12'h898;
    assign memory[7240] = 12'h898;
    assign memory[7241] = 12'h898;
    assign memory[7242] = 12'h898;
    assign memory[7243] = 12'h898;
    assign memory[7244] = 12'h898;
    assign memory[7245] = 12'h898;
    assign memory[7246] = 12'h898;
    assign memory[7247] = 12'h898;
    assign memory[7248] = 12'h898;
    assign memory[7249] = 12'h898;
    assign memory[7250] = 12'h898;
    assign memory[7251] = 12'h898;
    assign memory[7252] = 12'h898;
    assign memory[7253] = 12'h898;
    assign memory[7254] = 12'h898;
    assign memory[7255] = 12'h898;
    assign memory[7256] = 12'h898;
    assign memory[7257] = 12'h898;
    assign memory[7258] = 12'h898;
    assign memory[7259] = 12'h898;
    assign memory[7260] = 12'h898;
    assign memory[7261] = 12'h898;
    assign memory[7262] = 12'h898;
    assign memory[7263] = 12'h654;
    assign memory[7264] = 12'h654;
    assign memory[7265] = 12'h898;
    assign memory[7266] = 12'h898;
    assign memory[7267] = 12'hcbb;
    assign memory[7268] = 12'hcbb;
    assign memory[7269] = 12'hcbb;
    assign memory[7270] = 12'h898;
    assign memory[7271] = 12'h898;
    assign memory[7272] = 12'h898;
    assign memory[7273] = 12'h898;
    assign memory[7274] = 12'hcbb;
    assign memory[7275] = 12'hcbb;
    assign memory[7276] = 12'hcbb;
    assign memory[7277] = 12'hcbb;
    assign memory[7278] = 12'hcbb;
    assign memory[7279] = 12'hcbb;
    assign memory[7280] = 12'hcbb;
    assign memory[7281] = 12'hcbb;
    assign memory[7282] = 12'hcbb;
    assign memory[7283] = 12'h898;
    assign memory[7284] = 12'h898;
    assign memory[7285] = 12'h898;
    assign memory[7286] = 12'h898;
    assign memory[7287] = 12'h898;
    assign memory[7288] = 12'hcbb;
    assign memory[7289] = 12'hcbb;
    assign memory[7290] = 12'hcbb;
    assign memory[7291] = 12'hcbb;
    assign memory[7292] = 12'hcbb;
    assign memory[7293] = 12'h898;
    assign memory[7294] = 12'h898;
    assign memory[7295] = 12'h654;
    assign memory[7296] = 12'h654;
    assign memory[7297] = 12'h898;
    assign memory[7298] = 12'h898;
    assign memory[7299] = 12'hcbb;
    assign memory[7300] = 12'hcbb;
    assign memory[7301] = 12'hcbb;
    assign memory[7302] = 12'hcbb;
    assign memory[7303] = 12'hcbb;
    assign memory[7304] = 12'hcbb;
    assign memory[7305] = 12'hcbb;
    assign memory[7306] = 12'hcbb;
    assign memory[7307] = 12'hcbb;
    assign memory[7308] = 12'hcbb;
    assign memory[7309] = 12'hcbb;
    assign memory[7310] = 12'hcbb;
    assign memory[7311] = 12'hcbb;
    assign memory[7312] = 12'hcbb;
    assign memory[7313] = 12'hcbb;
    assign memory[7314] = 12'hcbb;
    assign memory[7315] = 12'hcbb;
    assign memory[7316] = 12'hcbb;
    assign memory[7317] = 12'hcbb;
    assign memory[7318] = 12'hcbb;
    assign memory[7319] = 12'hcbb;
    assign memory[7320] = 12'hcbb;
    assign memory[7321] = 12'hcbb;
    assign memory[7322] = 12'hcbb;
    assign memory[7323] = 12'hcbb;
    assign memory[7324] = 12'hcbb;
    assign memory[7325] = 12'h898;
    assign memory[7326] = 12'h898;
    assign memory[7327] = 12'h654;
    assign memory[7328] = 12'h654;
    assign memory[7329] = 12'h898;
    assign memory[7330] = 12'h898;
    assign memory[7331] = 12'hcbb;
    assign memory[7332] = 12'hcbb;
    assign memory[7333] = 12'hcbb;
    assign memory[7334] = 12'hcbb;
    assign memory[7335] = 12'hcbb;
    assign memory[7336] = 12'hcbb;
    assign memory[7337] = 12'hcbb;
    assign memory[7338] = 12'hcbb;
    assign memory[7339] = 12'hcbb;
    assign memory[7340] = 12'hcbb;
    assign memory[7341] = 12'hcbb;
    assign memory[7342] = 12'hcbb;
    assign memory[7343] = 12'hcbb;
    assign memory[7344] = 12'hcbb;
    assign memory[7345] = 12'hcbb;
    assign memory[7346] = 12'hcbb;
    assign memory[7347] = 12'hcbb;
    assign memory[7348] = 12'hcbb;
    assign memory[7349] = 12'hcbb;
    assign memory[7350] = 12'hcbb;
    assign memory[7351] = 12'hcbb;
    assign memory[7352] = 12'hcbb;
    assign memory[7353] = 12'haba;
    assign memory[7354] = 12'hcbb;
    assign memory[7355] = 12'hcbb;
    assign memory[7356] = 12'hcbb;
    assign memory[7357] = 12'h898;
    assign memory[7358] = 12'h898;
    assign memory[7359] = 12'h654;
    assign memory[7360] = 12'h654;
    assign memory[7361] = 12'h898;
    assign memory[7362] = 12'h898;
    assign memory[7363] = 12'h898;
    assign memory[7364] = 12'hcbb;
    assign memory[7365] = 12'hcbb;
    assign memory[7366] = 12'hcbb;
    assign memory[7367] = 12'hcbb;
    assign memory[7368] = 12'hcbb;
    assign memory[7369] = 12'hcbb;
    assign memory[7370] = 12'hcbb;
    assign memory[7371] = 12'hcbb;
    assign memory[7372] = 12'hcbb;
    assign memory[7373] = 12'hcbb;
    assign memory[7374] = 12'hcbb;
    assign memory[7375] = 12'hcbb;
    assign memory[7376] = 12'hcbb;
    assign memory[7377] = 12'hcbb;
    assign memory[7378] = 12'hcbb;
    assign memory[7379] = 12'hcbb;
    assign memory[7380] = 12'hcbb;
    assign memory[7381] = 12'hcbb;
    assign memory[7382] = 12'hcbb;
    assign memory[7383] = 12'hcbb;
    assign memory[7384] = 12'hcbb;
    assign memory[7385] = 12'hcbb;
    assign memory[7386] = 12'hcbb;
    assign memory[7387] = 12'hcbb;
    assign memory[7388] = 12'hcbb;
    assign memory[7389] = 12'h898;
    assign memory[7390] = 12'h898;
    assign memory[7391] = 12'h654;
    assign memory[7392] = 12'h654;
    assign memory[7393] = 12'h898;
    assign memory[7394] = 12'h898;
    assign memory[7395] = 12'h898;
    assign memory[7396] = 12'hcbb;
    assign memory[7397] = 12'hcbb;
    assign memory[7398] = 12'hcbb;
    assign memory[7399] = 12'hcbb;
    assign memory[7400] = 12'hcbb;
    assign memory[7401] = 12'hcbb;
    assign memory[7402] = 12'haba;
    assign memory[7403] = 12'hcbb;
    assign memory[7404] = 12'hcbb;
    assign memory[7405] = 12'hcbb;
    assign memory[7406] = 12'hcbb;
    assign memory[7407] = 12'hcbb;
    assign memory[7408] = 12'hcbb;
    assign memory[7409] = 12'hcbb;
    assign memory[7410] = 12'hcbb;
    assign memory[7411] = 12'hcbb;
    assign memory[7412] = 12'hcbb;
    assign memory[7413] = 12'hcbb;
    assign memory[7414] = 12'hcbb;
    assign memory[7415] = 12'hcbb;
    assign memory[7416] = 12'hcbb;
    assign memory[7417] = 12'hcbb;
    assign memory[7418] = 12'hcbb;
    assign memory[7419] = 12'hcbb;
    assign memory[7420] = 12'hcbb;
    assign memory[7421] = 12'h898;
    assign memory[7422] = 12'h898;
    assign memory[7423] = 12'h654;
    assign memory[7424] = 12'h654;
    assign memory[7425] = 12'h898;
    assign memory[7426] = 12'h898;
    assign memory[7427] = 12'h898;
    assign memory[7428] = 12'hcbb;
    assign memory[7429] = 12'hcbb;
    assign memory[7430] = 12'hcbb;
    assign memory[7431] = 12'hcbb;
    assign memory[7432] = 12'hcbb;
    assign memory[7433] = 12'hcbb;
    assign memory[7434] = 12'hcbb;
    assign memory[7435] = 12'hcbb;
    assign memory[7436] = 12'hcbb;
    assign memory[7437] = 12'hcbb;
    assign memory[7438] = 12'hcbb;
    assign memory[7439] = 12'hcbb;
    assign memory[7440] = 12'hcbb;
    assign memory[7441] = 12'hcbb;
    assign memory[7442] = 12'hcbb;
    assign memory[7443] = 12'hcbb;
    assign memory[7444] = 12'haba;
    assign memory[7445] = 12'hcbb;
    assign memory[7446] = 12'hcbb;
    assign memory[7447] = 12'hcbb;
    assign memory[7448] = 12'hcbb;
    assign memory[7449] = 12'hcbb;
    assign memory[7450] = 12'hcbb;
    assign memory[7451] = 12'hcbb;
    assign memory[7452] = 12'hcbb;
    assign memory[7453] = 12'h898;
    assign memory[7454] = 12'h898;
    assign memory[7455] = 12'h654;
    assign memory[7456] = 12'h654;
    assign memory[7457] = 12'h898;
    assign memory[7458] = 12'h898;
    assign memory[7459] = 12'hcbb;
    assign memory[7460] = 12'hcbb;
    assign memory[7461] = 12'hcbb;
    assign memory[7462] = 12'hcbb;
    assign memory[7463] = 12'hcbb;
    assign memory[7464] = 12'hcbb;
    assign memory[7465] = 12'hcbb;
    assign memory[7466] = 12'hcbb;
    assign memory[7467] = 12'hcbb;
    assign memory[7468] = 12'hcbb;
    assign memory[7469] = 12'hcbb;
    assign memory[7470] = 12'hcbb;
    assign memory[7471] = 12'hcbb;
    assign memory[7472] = 12'hcbb;
    assign memory[7473] = 12'hcbb;
    assign memory[7474] = 12'hcbb;
    assign memory[7475] = 12'hcbb;
    assign memory[7476] = 12'hcbb;
    assign memory[7477] = 12'hcbb;
    assign memory[7478] = 12'hcbb;
    assign memory[7479] = 12'hcbb;
    assign memory[7480] = 12'hcbb;
    assign memory[7481] = 12'hcbb;
    assign memory[7482] = 12'hcbb;
    assign memory[7483] = 12'hcbb;
    assign memory[7484] = 12'h898;
    assign memory[7485] = 12'h898;
    assign memory[7486] = 12'h898;
    assign memory[7487] = 12'h654;
    assign memory[7488] = 12'h654;
    assign memory[7489] = 12'h898;
    assign memory[7490] = 12'h898;
    assign memory[7491] = 12'hcbb;
    assign memory[7492] = 12'hcbb;
    assign memory[7493] = 12'hcbb;
    assign memory[7494] = 12'hcbb;
    assign memory[7495] = 12'hcbb;
    assign memory[7496] = 12'hcbb;
    assign memory[7497] = 12'hcbb;
    assign memory[7498] = 12'hcbb;
    assign memory[7499] = 12'hcbb;
    assign memory[7500] = 12'hcbb;
    assign memory[7501] = 12'hcbb;
    assign memory[7502] = 12'hcbb;
    assign memory[7503] = 12'hcbb;
    assign memory[7504] = 12'hcbb;
    assign memory[7505] = 12'hcbb;
    assign memory[7506] = 12'hcbb;
    assign memory[7507] = 12'hcbb;
    assign memory[7508] = 12'hcbb;
    assign memory[7509] = 12'hcbb;
    assign memory[7510] = 12'hcbb;
    assign memory[7511] = 12'hcbb;
    assign memory[7512] = 12'hcbb;
    assign memory[7513] = 12'hcbb;
    assign memory[7514] = 12'hcbb;
    assign memory[7515] = 12'hcbb;
    assign memory[7516] = 12'h898;
    assign memory[7517] = 12'h898;
    assign memory[7518] = 12'h898;
    assign memory[7519] = 12'h654;
    assign memory[7520] = 12'h654;
    assign memory[7521] = 12'h898;
    assign memory[7522] = 12'h898;
    assign memory[7523] = 12'hcbb;
    assign memory[7524] = 12'hcbb;
    assign memory[7525] = 12'hcbb;
    assign memory[7526] = 12'hcbb;
    assign memory[7527] = 12'hcbb;
    assign memory[7528] = 12'hcbb;
    assign memory[7529] = 12'hcbb;
    assign memory[7530] = 12'hcbb;
    assign memory[7531] = 12'hcbb;
    assign memory[7532] = 12'hcbb;
    assign memory[7533] = 12'hcbb;
    assign memory[7534] = 12'hcbb;
    assign memory[7535] = 12'haba;
    assign memory[7536] = 12'hcbb;
    assign memory[7537] = 12'hcbb;
    assign memory[7538] = 12'hcbb;
    assign memory[7539] = 12'hcbb;
    assign memory[7540] = 12'hcbb;
    assign memory[7541] = 12'hcbb;
    assign memory[7542] = 12'hcbb;
    assign memory[7543] = 12'hcbb;
    assign memory[7544] = 12'hcbb;
    assign memory[7545] = 12'hcbb;
    assign memory[7546] = 12'hcbb;
    assign memory[7547] = 12'hcbb;
    assign memory[7548] = 12'h898;
    assign memory[7549] = 12'h898;
    assign memory[7550] = 12'h898;
    assign memory[7551] = 12'h654;
    assign memory[7552] = 12'h654;
    assign memory[7553] = 12'h898;
    assign memory[7554] = 12'h898;
    assign memory[7555] = 12'hcbb;
    assign memory[7556] = 12'hcbb;
    assign memory[7557] = 12'hcbb;
    assign memory[7558] = 12'hcbb;
    assign memory[7559] = 12'hcbb;
    assign memory[7560] = 12'hcbb;
    assign memory[7561] = 12'hcbb;
    assign memory[7562] = 12'hcbb;
    assign memory[7563] = 12'hcbb;
    assign memory[7564] = 12'hcbb;
    assign memory[7565] = 12'hcbb;
    assign memory[7566] = 12'hcbb;
    assign memory[7567] = 12'hcbb;
    assign memory[7568] = 12'hcbb;
    assign memory[7569] = 12'hcbb;
    assign memory[7570] = 12'hcbb;
    assign memory[7571] = 12'hcbb;
    assign memory[7572] = 12'hcbb;
    assign memory[7573] = 12'hcbb;
    assign memory[7574] = 12'hcbb;
    assign memory[7575] = 12'hcbb;
    assign memory[7576] = 12'hcbb;
    assign memory[7577] = 12'hcbb;
    assign memory[7578] = 12'hcbb;
    assign memory[7579] = 12'hcbb;
    assign memory[7580] = 12'h898;
    assign memory[7581] = 12'h898;
    assign memory[7582] = 12'h898;
    assign memory[7583] = 12'h654;
    assign memory[7584] = 12'h654;
    assign memory[7585] = 12'h898;
    assign memory[7586] = 12'h898;
    assign memory[7587] = 12'hcbb;
    assign memory[7588] = 12'hcbb;
    assign memory[7589] = 12'hcbb;
    assign memory[7590] = 12'hcbb;
    assign memory[7591] = 12'hcbb;
    assign memory[7592] = 12'hcbb;
    assign memory[7593] = 12'hcbb;
    assign memory[7594] = 12'hcbb;
    assign memory[7595] = 12'hcbb;
    assign memory[7596] = 12'hcbb;
    assign memory[7597] = 12'hcbb;
    assign memory[7598] = 12'hcbb;
    assign memory[7599] = 12'hcbb;
    assign memory[7600] = 12'hcbb;
    assign memory[7601] = 12'hcbb;
    assign memory[7602] = 12'hcbb;
    assign memory[7603] = 12'hcbb;
    assign memory[7604] = 12'hcbb;
    assign memory[7605] = 12'hcbb;
    assign memory[7606] = 12'hcbb;
    assign memory[7607] = 12'hcbb;
    assign memory[7608] = 12'hcbb;
    assign memory[7609] = 12'hcbb;
    assign memory[7610] = 12'hcbb;
    assign memory[7611] = 12'hcbb;
    assign memory[7612] = 12'h898;
    assign memory[7613] = 12'h898;
    assign memory[7614] = 12'h898;
    assign memory[7615] = 12'h654;
    assign memory[7616] = 12'h654;
    assign memory[7617] = 12'h898;
    assign memory[7618] = 12'h898;
    assign memory[7619] = 12'hcbb;
    assign memory[7620] = 12'hcbb;
    assign memory[7621] = 12'hcbb;
    assign memory[7622] = 12'hcbb;
    assign memory[7623] = 12'hcbb;
    assign memory[7624] = 12'haba;
    assign memory[7625] = 12'hcbb;
    assign memory[7626] = 12'hcbb;
    assign memory[7627] = 12'hcbb;
    assign memory[7628] = 12'hcbb;
    assign memory[7629] = 12'hcbb;
    assign memory[7630] = 12'haba;
    assign memory[7631] = 12'hcbb;
    assign memory[7632] = 12'hcbb;
    assign memory[7633] = 12'hcbb;
    assign memory[7634] = 12'hcbb;
    assign memory[7635] = 12'hcbb;
    assign memory[7636] = 12'hcbb;
    assign memory[7637] = 12'hcbb;
    assign memory[7638] = 12'haba;
    assign memory[7639] = 12'hcbb;
    assign memory[7640] = 12'hcbb;
    assign memory[7641] = 12'hcbb;
    assign memory[7642] = 12'hcbb;
    assign memory[7643] = 12'hcbb;
    assign memory[7644] = 12'hcbb;
    assign memory[7645] = 12'h898;
    assign memory[7646] = 12'h898;
    assign memory[7647] = 12'h654;
    assign memory[7648] = 12'h654;
    assign memory[7649] = 12'h898;
    assign memory[7650] = 12'h898;
    assign memory[7651] = 12'hcbb;
    assign memory[7652] = 12'hcbb;
    assign memory[7653] = 12'hcbb;
    assign memory[7654] = 12'hcbb;
    assign memory[7655] = 12'hcbb;
    assign memory[7656] = 12'hcbb;
    assign memory[7657] = 12'hcbb;
    assign memory[7658] = 12'hcbb;
    assign memory[7659] = 12'hcbb;
    assign memory[7660] = 12'hcbb;
    assign memory[7661] = 12'hcbb;
    assign memory[7662] = 12'hcbb;
    assign memory[7663] = 12'hcbb;
    assign memory[7664] = 12'hcbb;
    assign memory[7665] = 12'hcbb;
    assign memory[7666] = 12'hcbb;
    assign memory[7667] = 12'hcbb;
    assign memory[7668] = 12'hcbb;
    assign memory[7669] = 12'hcbb;
    assign memory[7670] = 12'hcbb;
    assign memory[7671] = 12'hcbb;
    assign memory[7672] = 12'hcbb;
    assign memory[7673] = 12'hcbb;
    assign memory[7674] = 12'hcbb;
    assign memory[7675] = 12'hcbb;
    assign memory[7676] = 12'hcbb;
    assign memory[7677] = 12'h898;
    assign memory[7678] = 12'h898;
    assign memory[7679] = 12'h654;
    assign memory[7680] = 12'h654;
    assign memory[7681] = 12'h898;
    assign memory[7682] = 12'h898;
    assign memory[7683] = 12'hcbb;
    assign memory[7684] = 12'hcbb;
    assign memory[7685] = 12'hcbb;
    assign memory[7686] = 12'hcbb;
    assign memory[7687] = 12'hcbb;
    assign memory[7688] = 12'hcbb;
    assign memory[7689] = 12'hcbb;
    assign memory[7690] = 12'hcbb;
    assign memory[7691] = 12'hcbb;
    assign memory[7692] = 12'hcbb;
    assign memory[7693] = 12'hcbb;
    assign memory[7694] = 12'hcbb;
    assign memory[7695] = 12'hcbb;
    assign memory[7696] = 12'hcbb;
    assign memory[7697] = 12'hcbb;
    assign memory[7698] = 12'hcbb;
    assign memory[7699] = 12'hcbb;
    assign memory[7700] = 12'hcbb;
    assign memory[7701] = 12'hcbb;
    assign memory[7702] = 12'hcbb;
    assign memory[7703] = 12'hcbb;
    assign memory[7704] = 12'hcbb;
    assign memory[7705] = 12'hcbb;
    assign memory[7706] = 12'hcbb;
    assign memory[7707] = 12'hcbb;
    assign memory[7708] = 12'hcbb;
    assign memory[7709] = 12'h898;
    assign memory[7710] = 12'h898;
    assign memory[7711] = 12'h654;
    assign memory[7712] = 12'h654;
    assign memory[7713] = 12'h898;
    assign memory[7714] = 12'h898;
    assign memory[7715] = 12'hcbb;
    assign memory[7716] = 12'hcbb;
    assign memory[7717] = 12'hcbb;
    assign memory[7718] = 12'hcbb;
    assign memory[7719] = 12'hcbb;
    assign memory[7720] = 12'hcbb;
    assign memory[7721] = 12'hcbb;
    assign memory[7722] = 12'hcbb;
    assign memory[7723] = 12'hcbb;
    assign memory[7724] = 12'hcbb;
    assign memory[7725] = 12'hcbb;
    assign memory[7726] = 12'hcbb;
    assign memory[7727] = 12'hcbb;
    assign memory[7728] = 12'haba;
    assign memory[7729] = 12'hcbb;
    assign memory[7730] = 12'hcbb;
    assign memory[7731] = 12'hcbb;
    assign memory[7732] = 12'hcbb;
    assign memory[7733] = 12'hcbb;
    assign memory[7734] = 12'hcbb;
    assign memory[7735] = 12'hcbb;
    assign memory[7736] = 12'hcbb;
    assign memory[7737] = 12'hcbb;
    assign memory[7738] = 12'hcbb;
    assign memory[7739] = 12'hcbb;
    assign memory[7740] = 12'hcbb;
    assign memory[7741] = 12'h898;
    assign memory[7742] = 12'h898;
    assign memory[7743] = 12'h654;
    assign memory[7744] = 12'h654;
    assign memory[7745] = 12'h898;
    assign memory[7746] = 12'h898;
    assign memory[7747] = 12'hcbb;
    assign memory[7748] = 12'hcbb;
    assign memory[7749] = 12'hcbb;
    assign memory[7750] = 12'hcbb;
    assign memory[7751] = 12'hcbb;
    assign memory[7752] = 12'hcbb;
    assign memory[7753] = 12'hcbb;
    assign memory[7754] = 12'hcbb;
    assign memory[7755] = 12'hcbb;
    assign memory[7756] = 12'hcbb;
    assign memory[7757] = 12'hcbb;
    assign memory[7758] = 12'hcbb;
    assign memory[7759] = 12'hcbb;
    assign memory[7760] = 12'hcbb;
    assign memory[7761] = 12'hcbb;
    assign memory[7762] = 12'hcbb;
    assign memory[7763] = 12'hcbb;
    assign memory[7764] = 12'hcbb;
    assign memory[7765] = 12'hcbb;
    assign memory[7766] = 12'hcbb;
    assign memory[7767] = 12'hcbb;
    assign memory[7768] = 12'hcbb;
    assign memory[7769] = 12'haba;
    assign memory[7770] = 12'hcbb;
    assign memory[7771] = 12'hcbb;
    assign memory[7772] = 12'h898;
    assign memory[7773] = 12'h898;
    assign memory[7774] = 12'h898;
    assign memory[7775] = 12'h654;
    assign memory[7776] = 12'h654;
    assign memory[7777] = 12'h898;
    assign memory[7778] = 12'h898;
    assign memory[7779] = 12'h898;
    assign memory[7780] = 12'hcbb;
    assign memory[7781] = 12'hcbb;
    assign memory[7782] = 12'hcbb;
    assign memory[7783] = 12'hcbb;
    assign memory[7784] = 12'hcbb;
    assign memory[7785] = 12'hcbb;
    assign memory[7786] = 12'hcbb;
    assign memory[7787] = 12'hcbb;
    assign memory[7788] = 12'hcbb;
    assign memory[7789] = 12'hcbb;
    assign memory[7790] = 12'hcbb;
    assign memory[7791] = 12'hcbb;
    assign memory[7792] = 12'hcbb;
    assign memory[7793] = 12'hcbb;
    assign memory[7794] = 12'hcbb;
    assign memory[7795] = 12'hcbb;
    assign memory[7796] = 12'hcbb;
    assign memory[7797] = 12'hcbb;
    assign memory[7798] = 12'hcbb;
    assign memory[7799] = 12'hcbb;
    assign memory[7800] = 12'hcbb;
    assign memory[7801] = 12'haba;
    assign memory[7802] = 12'hcbb;
    assign memory[7803] = 12'hcbb;
    assign memory[7804] = 12'h898;
    assign memory[7805] = 12'h898;
    assign memory[7806] = 12'h898;
    assign memory[7807] = 12'h654;
    assign memory[7808] = 12'h654;
    assign memory[7809] = 12'h898;
    assign memory[7810] = 12'h898;
    assign memory[7811] = 12'h898;
    assign memory[7812] = 12'hcbb;
    assign memory[7813] = 12'hcbb;
    assign memory[7814] = 12'hcbb;
    assign memory[7815] = 12'hcbb;
    assign memory[7816] = 12'hcbb;
    assign memory[7817] = 12'hcbb;
    assign memory[7818] = 12'hcbb;
    assign memory[7819] = 12'hcbb;
    assign memory[7820] = 12'hcbb;
    assign memory[7821] = 12'hcbb;
    assign memory[7822] = 12'hcbb;
    assign memory[7823] = 12'hcbb;
    assign memory[7824] = 12'hcbb;
    assign memory[7825] = 12'hcbb;
    assign memory[7826] = 12'hcbb;
    assign memory[7827] = 12'hcbb;
    assign memory[7828] = 12'hcbb;
    assign memory[7829] = 12'hcbb;
    assign memory[7830] = 12'hcbb;
    assign memory[7831] = 12'hcbb;
    assign memory[7832] = 12'hcbb;
    assign memory[7833] = 12'hcbb;
    assign memory[7834] = 12'hcbb;
    assign memory[7835] = 12'hcbb;
    assign memory[7836] = 12'h898;
    assign memory[7837] = 12'h898;
    assign memory[7838] = 12'h898;
    assign memory[7839] = 12'h654;
    assign memory[7840] = 12'h654;
    assign memory[7841] = 12'h898;
    assign memory[7842] = 12'h898;
    assign memory[7843] = 12'h898;
    assign memory[7844] = 12'hcbb;
    assign memory[7845] = 12'hcbb;
    assign memory[7846] = 12'hcbb;
    assign memory[7847] = 12'hcbb;
    assign memory[7848] = 12'hcbb;
    assign memory[7849] = 12'hcbb;
    assign memory[7850] = 12'hcbb;
    assign memory[7851] = 12'hcbb;
    assign memory[7852] = 12'hcbb;
    assign memory[7853] = 12'hcbb;
    assign memory[7854] = 12'hcbb;
    assign memory[7855] = 12'hcbb;
    assign memory[7856] = 12'hcbb;
    assign memory[7857] = 12'hcbb;
    assign memory[7858] = 12'hcbb;
    assign memory[7859] = 12'hcbb;
    assign memory[7860] = 12'hcbb;
    assign memory[7861] = 12'hcbb;
    assign memory[7862] = 12'hcbb;
    assign memory[7863] = 12'hcbb;
    assign memory[7864] = 12'hcbb;
    assign memory[7865] = 12'hcbb;
    assign memory[7866] = 12'hcbb;
    assign memory[7867] = 12'hcbb;
    assign memory[7868] = 12'h898;
    assign memory[7869] = 12'h898;
    assign memory[7870] = 12'h898;
    assign memory[7871] = 12'h654;
    assign memory[7872] = 12'h654;
    assign memory[7873] = 12'h898;
    assign memory[7874] = 12'h898;
    assign memory[7875] = 12'h898;
    assign memory[7876] = 12'hcbb;
    assign memory[7877] = 12'hcbb;
    assign memory[7878] = 12'hcbb;
    assign memory[7879] = 12'hcbb;
    assign memory[7880] = 12'hcbb;
    assign memory[7881] = 12'hcbb;
    assign memory[7882] = 12'hcbb;
    assign memory[7883] = 12'hcbb;
    assign memory[7884] = 12'hcbb;
    assign memory[7885] = 12'haba;
    assign memory[7886] = 12'hcbb;
    assign memory[7887] = 12'hcbb;
    assign memory[7888] = 12'hcbb;
    assign memory[7889] = 12'hcbb;
    assign memory[7890] = 12'hcbb;
    assign memory[7891] = 12'hcbb;
    assign memory[7892] = 12'hcbb;
    assign memory[7893] = 12'hcbb;
    assign memory[7894] = 12'hcbb;
    assign memory[7895] = 12'hcbb;
    assign memory[7896] = 12'hcbb;
    assign memory[7897] = 12'hcbb;
    assign memory[7898] = 12'hcbb;
    assign memory[7899] = 12'hcbb;
    assign memory[7900] = 12'hcbb;
    assign memory[7901] = 12'h898;
    assign memory[7902] = 12'h898;
    assign memory[7903] = 12'h654;
    assign memory[7904] = 12'h654;
    assign memory[7905] = 12'h898;
    assign memory[7906] = 12'h898;
    assign memory[7907] = 12'h898;
    assign memory[7908] = 12'hcbb;
    assign memory[7909] = 12'hcbb;
    assign memory[7910] = 12'hcbb;
    assign memory[7911] = 12'hcbb;
    assign memory[7912] = 12'haba;
    assign memory[7913] = 12'hcbb;
    assign memory[7914] = 12'hcbb;
    assign memory[7915] = 12'hcbb;
    assign memory[7916] = 12'hcbb;
    assign memory[7917] = 12'hcbb;
    assign memory[7918] = 12'hcbb;
    assign memory[7919] = 12'hcbb;
    assign memory[7920] = 12'hcbb;
    assign memory[7921] = 12'hcbb;
    assign memory[7922] = 12'hcbb;
    assign memory[7923] = 12'hcbb;
    assign memory[7924] = 12'hcbb;
    assign memory[7925] = 12'hcbb;
    assign memory[7926] = 12'haba;
    assign memory[7927] = 12'hcbb;
    assign memory[7928] = 12'hcbb;
    assign memory[7929] = 12'hcbb;
    assign memory[7930] = 12'hcbb;
    assign memory[7931] = 12'hcbb;
    assign memory[7932] = 12'hcbb;
    assign memory[7933] = 12'h898;
    assign memory[7934] = 12'h898;
    assign memory[7935] = 12'h654;
    assign memory[7936] = 12'h654;
    assign memory[7937] = 12'h898;
    assign memory[7938] = 12'h898;
    assign memory[7939] = 12'hcbb;
    assign memory[7940] = 12'hcbb;
    assign memory[7941] = 12'hcbb;
    assign memory[7942] = 12'hcbb;
    assign memory[7943] = 12'hcbb;
    assign memory[7944] = 12'hcbb;
    assign memory[7945] = 12'hcbb;
    assign memory[7946] = 12'hcbb;
    assign memory[7947] = 12'hcbb;
    assign memory[7948] = 12'hcbb;
    assign memory[7949] = 12'hcbb;
    assign memory[7950] = 12'hcbb;
    assign memory[7951] = 12'hcbb;
    assign memory[7952] = 12'hcbb;
    assign memory[7953] = 12'hcbb;
    assign memory[7954] = 12'hcbb;
    assign memory[7955] = 12'hcbb;
    assign memory[7956] = 12'hcbb;
    assign memory[7957] = 12'hcbb;
    assign memory[7958] = 12'hcbb;
    assign memory[7959] = 12'hcbb;
    assign memory[7960] = 12'hcbb;
    assign memory[7961] = 12'hcbb;
    assign memory[7962] = 12'hcbb;
    assign memory[7963] = 12'hcbb;
    assign memory[7964] = 12'hcbb;
    assign memory[7965] = 12'h898;
    assign memory[7966] = 12'h898;
    assign memory[7967] = 12'h654;
    assign memory[7968] = 12'h654;
    assign memory[7969] = 12'h898;
    assign memory[7970] = 12'h898;
    assign memory[7971] = 12'hcbb;
    assign memory[7972] = 12'hcbb;
    assign memory[7973] = 12'hcbb;
    assign memory[7974] = 12'hcbb;
    assign memory[7975] = 12'hcbb;
    assign memory[7976] = 12'hcbb;
    assign memory[7977] = 12'hcbb;
    assign memory[7978] = 12'hcbb;
    assign memory[7979] = 12'hcbb;
    assign memory[7980] = 12'hcbb;
    assign memory[7981] = 12'hcbb;
    assign memory[7982] = 12'hcbb;
    assign memory[7983] = 12'hcbb;
    assign memory[7984] = 12'hcbb;
    assign memory[7985] = 12'hcbb;
    assign memory[7986] = 12'hcbb;
    assign memory[7987] = 12'hcbb;
    assign memory[7988] = 12'hcbb;
    assign memory[7989] = 12'hcbb;
    assign memory[7990] = 12'hcbb;
    assign memory[7991] = 12'hcbb;
    assign memory[7992] = 12'hcbb;
    assign memory[7993] = 12'hcbb;
    assign memory[7994] = 12'haba;
    assign memory[7995] = 12'hcbb;
    assign memory[7996] = 12'hcbb;
    assign memory[7997] = 12'h898;
    assign memory[7998] = 12'h898;
    assign memory[7999] = 12'h654;
    assign memory[8000] = 12'h654;
    assign memory[8001] = 12'h898;
    assign memory[8002] = 12'h898;
    assign memory[8003] = 12'hcbb;
    assign memory[8004] = 12'hcbb;
    assign memory[8005] = 12'hcbb;
    assign memory[8006] = 12'hcbb;
    assign memory[8007] = 12'hcbb;
    assign memory[8008] = 12'hcbb;
    assign memory[8009] = 12'hcbb;
    assign memory[8010] = 12'hcbb;
    assign memory[8011] = 12'hcbb;
    assign memory[8012] = 12'hcbb;
    assign memory[8013] = 12'hcbb;
    assign memory[8014] = 12'hcbb;
    assign memory[8015] = 12'hcbb;
    assign memory[8016] = 12'hcbb;
    assign memory[8017] = 12'hcbb;
    assign memory[8018] = 12'hcbb;
    assign memory[8019] = 12'hcbb;
    assign memory[8020] = 12'hcbb;
    assign memory[8021] = 12'hcbb;
    assign memory[8022] = 12'hcbb;
    assign memory[8023] = 12'hcbb;
    assign memory[8024] = 12'hcbb;
    assign memory[8025] = 12'hcbb;
    assign memory[8026] = 12'hcbb;
    assign memory[8027] = 12'hcbb;
    assign memory[8028] = 12'h898;
    assign memory[8029] = 12'h898;
    assign memory[8030] = 12'h898;
    assign memory[8031] = 12'h654;
    assign memory[8032] = 12'h654;
    assign memory[8033] = 12'h898;
    assign memory[8034] = 12'h898;
    assign memory[8035] = 12'hcbb;
    assign memory[8036] = 12'hcbb;
    assign memory[8037] = 12'hcbb;
    assign memory[8038] = 12'hcbb;
    assign memory[8039] = 12'hcbb;
    assign memory[8040] = 12'hcbb;
    assign memory[8041] = 12'hcbb;
    assign memory[8042] = 12'hcbb;
    assign memory[8043] = 12'hcbb;
    assign memory[8044] = 12'hcbb;
    assign memory[8045] = 12'hcbb;
    assign memory[8046] = 12'hcbb;
    assign memory[8047] = 12'hcbb;
    assign memory[8048] = 12'hcbb;
    assign memory[8049] = 12'hcbb;
    assign memory[8050] = 12'hcbb;
    assign memory[8051] = 12'hcbb;
    assign memory[8052] = 12'hcbb;
    assign memory[8053] = 12'hcbb;
    assign memory[8054] = 12'hcbb;
    assign memory[8055] = 12'hcbb;
    assign memory[8056] = 12'hcbb;
    assign memory[8057] = 12'hcbb;
    assign memory[8058] = 12'hcbb;
    assign memory[8059] = 12'hcbb;
    assign memory[8060] = 12'h898;
    assign memory[8061] = 12'h898;
    assign memory[8062] = 12'h898;
    assign memory[8063] = 12'h654;
    assign memory[8064] = 12'h654;
    assign memory[8065] = 12'h898;
    assign memory[8066] = 12'h898;
    assign memory[8067] = 12'hcbb;
    assign memory[8068] = 12'hcbb;
    assign memory[8069] = 12'hcbb;
    assign memory[8070] = 12'hcbb;
    assign memory[8071] = 12'h898;
    assign memory[8072] = 12'h898;
    assign memory[8073] = 12'h898;
    assign memory[8074] = 12'h898;
    assign memory[8075] = 12'hcbb;
    assign memory[8076] = 12'hcbb;
    assign memory[8077] = 12'hcbb;
    assign memory[8078] = 12'h898;
    assign memory[8079] = 12'h898;
    assign memory[8080] = 12'h898;
    assign memory[8081] = 12'hcbb;
    assign memory[8082] = 12'hcbb;
    assign memory[8083] = 12'hcbb;
    assign memory[8084] = 12'hcbb;
    assign memory[8085] = 12'h898;
    assign memory[8086] = 12'h898;
    assign memory[8087] = 12'h898;
    assign memory[8088] = 12'hcbb;
    assign memory[8089] = 12'hcbb;
    assign memory[8090] = 12'hcbb;
    assign memory[8091] = 12'hcbb;
    assign memory[8092] = 12'hcbb;
    assign memory[8093] = 12'h898;
    assign memory[8094] = 12'h898;
    assign memory[8095] = 12'h654;
    assign memory[8096] = 12'h654;
    assign memory[8097] = 12'h898;
    assign memory[8098] = 12'h898;
    assign memory[8099] = 12'h898;
    assign memory[8100] = 12'h898;
    assign memory[8101] = 12'h898;
    assign memory[8102] = 12'h898;
    assign memory[8103] = 12'h898;
    assign memory[8104] = 12'h898;
    assign memory[8105] = 12'h898;
    assign memory[8106] = 12'h898;
    assign memory[8107] = 12'h898;
    assign memory[8108] = 12'h898;
    assign memory[8109] = 12'h898;
    assign memory[8110] = 12'h898;
    assign memory[8111] = 12'h898;
    assign memory[8112] = 12'h898;
    assign memory[8113] = 12'h898;
    assign memory[8114] = 12'h898;
    assign memory[8115] = 12'h898;
    assign memory[8116] = 12'h898;
    assign memory[8117] = 12'h898;
    assign memory[8118] = 12'h898;
    assign memory[8119] = 12'h898;
    assign memory[8120] = 12'h898;
    assign memory[8121] = 12'h898;
    assign memory[8122] = 12'h898;
    assign memory[8123] = 12'h898;
    assign memory[8124] = 12'h898;
    assign memory[8125] = 12'h898;
    assign memory[8126] = 12'h898;
    assign memory[8127] = 12'h654;
    assign memory[8128] = 12'h654;
    assign memory[8129] = 12'h898;
    assign memory[8130] = 12'h898;
    assign memory[8131] = 12'h898;
    assign memory[8132] = 12'h898;
    assign memory[8133] = 12'h898;
    assign memory[8134] = 12'h898;
    assign memory[8135] = 12'h898;
    assign memory[8136] = 12'h898;
    assign memory[8137] = 12'h898;
    assign memory[8138] = 12'h898;
    assign memory[8139] = 12'h898;
    assign memory[8140] = 12'h898;
    assign memory[8141] = 12'h898;
    assign memory[8142] = 12'h898;
    assign memory[8143] = 12'h898;
    assign memory[8144] = 12'h898;
    assign memory[8145] = 12'h898;
    assign memory[8146] = 12'h898;
    assign memory[8147] = 12'h898;
    assign memory[8148] = 12'h898;
    assign memory[8149] = 12'h898;
    assign memory[8150] = 12'h898;
    assign memory[8151] = 12'h898;
    assign memory[8152] = 12'h898;
    assign memory[8153] = 12'h898;
    assign memory[8154] = 12'h898;
    assign memory[8155] = 12'h898;
    assign memory[8156] = 12'h898;
    assign memory[8157] = 12'h898;
    assign memory[8158] = 12'h898;
    assign memory[8159] = 12'h654;
    assign memory[8160] = 12'h654;
    assign memory[8161] = 12'h654;
    assign memory[8162] = 12'h654;
    assign memory[8163] = 12'h654;
    assign memory[8164] = 12'h654;
    assign memory[8165] = 12'h654;
    assign memory[8166] = 12'h654;
    assign memory[8167] = 12'h654;
    assign memory[8168] = 12'h654;
    assign memory[8169] = 12'h654;
    assign memory[8170] = 12'h654;
    assign memory[8171] = 12'h654;
    assign memory[8172] = 12'h654;
    assign memory[8173] = 12'h654;
    assign memory[8174] = 12'h654;
    assign memory[8175] = 12'h654;
    assign memory[8176] = 12'h654;
    assign memory[8177] = 12'h654;
    assign memory[8178] = 12'h654;
    assign memory[8179] = 12'h654;
    assign memory[8180] = 12'h654;
    assign memory[8181] = 12'h654;
    assign memory[8182] = 12'h654;
    assign memory[8183] = 12'h654;
    assign memory[8184] = 12'h654;
    assign memory[8185] = 12'h654;
    assign memory[8186] = 12'h654;
    assign memory[8187] = 12'h654;
    assign memory[8188] = 12'h654;
    assign memory[8189] = 12'h654;
    assign memory[8190] = 12'h654;
    assign memory[8191] = 12'h654;
endmodule