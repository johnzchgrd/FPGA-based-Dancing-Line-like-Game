//	How to use:	
//	1. Edit the songs on the Enter Song sheet.	
// 	2. Select this whole worksheet, copy it, and paste it into a new file.	
//	3. Save the file as song_rom.v.	

module saw2_rom (
    input clk,						
	output reg [25:0] dout,						
	input [11:0] addr		
    );
        
    wire [25:0] memory [4095:0];  			
	always @(posedge clk)						
		dout = memory[addr];					

    parameter s1 = 142;
    parameter s2 = s1 + 140;
    parameter s3 = s2 + 81;

    assign memory[0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[79 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[80 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[81 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[82 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[83 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[84 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[85 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[86 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[87 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[88 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[89 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[90 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[91 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[92 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[93 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[94 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[95 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[96 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[97 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[98 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[99 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[100] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[101] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[102] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[103] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[104] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[105] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[106] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[107] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[108] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[109] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[110] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[111] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[112] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[113] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[114] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[115] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[116] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[117] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[118] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[119] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[120] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[121] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[122] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[123] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[124] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[125] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[126] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[127] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[128] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[129] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[130] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[131] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[132] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[133] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[134] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[135] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[136] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[137] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[138] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[139] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[140] = {7'd0  , 8'd123, 7'd0  , 2'd0, 2'd0};
    assign memory[141] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s1+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s1+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+25 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+26 ] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+27 ] = {7'd31 , 8'd81 , 7'd112, 2'd0, 2'd0};
    assign memory[s1+28 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+29 ] = {7'd31 , 8'd24 , 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+30 ] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+31 ] = {7'd31 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+32 ] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+33 ] = {7'd31 , 8'd81 , 7'd112, 2'd0, 2'd0};
    assign memory[s1+34 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+35 ] = {7'd31 , 8'd24 , 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+36 ] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+37 ] = {7'd31 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+38 ] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+39 ] = {7'd31 , 8'd81 , 7'd112, 2'd0, 2'd0};
    assign memory[s1+40 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+41 ] = {7'd31 , 8'd24 , 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+42 ] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+43 ] = {7'd31 , 8'd129, 7'd112, 2'd0, 2'd0};
    assign memory[s1+44 ] = {7'd31 , 8'd255, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+45 ] = {7'd31 , 8'd81 , 7'd112, 2'd0, 2'd0};
    assign memory[s1+46 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+47 ] = {7'd31 , 8'd24 , 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+48 ] = {7'd31 , 8'd192, 7'd112, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+49 ] = {7'd27 , 8'd32 , 7'd112, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+50 ] = {7'd0  , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+51 ] = {7'd27 , 8'd32 , 7'd112, 2'd0, 2'd0};   //note: 3B
    assign memory[s1+52 ] = {7'd29 , 8'd32 , 7'd112, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+53 ] = {7'd0  , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+54 ] = {7'd29 , 8'd32 , 7'd112, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s1+55 ] = {7'd31 , 8'd72 , 7'd114, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s1+56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+79 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+80 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+81 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+82 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+83 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+84 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+85 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+86 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+87 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+88 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+89 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+90 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+91 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+92 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+93 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+94 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+95 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+96 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+97 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+98 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+99 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+100] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+101] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+102] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+103] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+104] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+105] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+106] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+107] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+108] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+109] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+110] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+111] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+112] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+113] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+114] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+115] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+116] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+117] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+118] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+119] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+120] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+121] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+122] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+123] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+124] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+125] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+126] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+127] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+128] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+129] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+130] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+131] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+132] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+133] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+134] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+135] = {7'd0  , 8'd135, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+136] = {7'd0  , 8'd1  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+137] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+138] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+139] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s2+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s2+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+79 ] = {7'd0  , 8'd79 , 7'd0  , 2'd0, 2'd0};
    assign memory[s2+80 ] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s3+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s3+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+74 ] = {7'd0  , 8'd107, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+75 ] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

endmodule							
