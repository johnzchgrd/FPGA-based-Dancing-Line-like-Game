`timescale 1ns / 1ps

module turn_points_rom(
    input                   clk,
    input                   reset,
    input                   load_raw,
    input [ 1:0]            song,
    input [10:0]            refer_x, refer_y,
    input [ 9:0]            current_block_x, current_block_y,
    input [ 9:0]            x1, y1, x2, y2,
    output reg              fail,
    output                  is_road,
    output [2:0]            debug
    );
 
    reg                     load;
    wire                    shift_enable;
    reg  [ 8:0]             cnt, cnt_next;
    wire [21:0]             memory  [453:0];
    wire [21:0]             memory2 [428:0];
    wire [21:0]             memory3 [186:0];
    wire [21:0]             memory4 [240:0];
    // turn point registers
    reg [21:0] turn1, turn2, turn3, turn4, turn5, turn6, turn7, turn8, turn9, 
				turn10, turn11, turn12, turn13, turn14, turn15, turn16, turn17, 
				turn18;
	wire scan_in_turn12, scan_in_turn23, scan_in_turn34, scan_in_turn45, scan_in_turn56, scan_in_turn67, scan_in_turn78, scan_in_turn89, scan_in_turn910, 
				scan_in_turn1011, scan_in_turn1112, scan_in_turn1213, scan_in_turn1314, scan_in_turn1415, scan_in_turn1516, scan_in_turn1617, scan_in_turn1718;
				
	wire dot1_in_turn12, dot1_in_turn23, dot1_in_turn34, dot1_in_turn45, dot1_in_turn56, dot1_in_turn67, dot1_in_turn78, dot1_in_turn89, dot1_in_turn910, 
				dot1_in_turn1011, dot1_in_turn1112, dot1_in_turn1213, dot1_in_turn1314, dot1_in_turn1415, dot1_in_turn1516, dot1_in_turn1617, dot1_in_turn1718;
				
	wire dot2_in_turn12, dot2_in_turn23, dot2_in_turn34, dot2_in_turn45, dot2_in_turn56, dot2_in_turn67, dot2_in_turn78, dot2_in_turn89, dot2_in_turn910, 
				dot2_in_turn1011, dot2_in_turn1112, dot2_in_turn1213, dot2_in_turn1314, dot2_in_turn1415, dot2_in_turn1516, dot2_in_turn1617, dot2_in_turn1718;
				
    //debug
    assign debug = {shift_enable,load_raw,fail}; 
    // judge when to update coordinate
    assign shift_enable = (turn2[21:11] <= refer_x + 21) & (turn2[10:0] <= refer_y + 16);
    //
    // ─── SHIFT REGISTER FILES ───────────────────────────────────────────────────────
    //

    always@(posedge clk) begin
        load <= load_raw;
        if(load) begin //initialize route
			case(song)
				2'd0: begin
					turn1 <= memory[16]; turn2 <= memory[15]; turn3 <= memory[14]; 
					turn4 <= memory[13]; turn5 <= memory[12]; turn6 <= memory[11]; 
					turn7 <= memory[10]; turn8 <= memory[ 9]; turn9 <= memory[ 8]; 
					turn10 <= memory[ 7]; turn11 <= memory[ 6]; turn12 <= memory[ 5]; 
					turn13 <= memory[ 4]; turn14 <= memory[ 3]; turn15 <= memory[ 2]; 
					turn16 <= memory[ 1]; turn17 <= memory[ 0]; turn18 <= memory[ 0]; 
				end
				2'd1: begin
					turn1 <= memory2[16]; turn2 <= memory2[15]; turn3 <= memory2[14]; 
					turn4 <= memory2[13]; turn5 <= memory2[12]; turn6 <= memory2[11]; 
					turn7 <= memory2[10]; turn8 <= memory2[ 9]; turn9 <= memory2[ 8]; 
					turn10 <= memory2[ 7]; turn11 <= memory2[ 6]; turn12 <= memory2[ 5]; 
					turn13 <= memory2[ 4]; turn14 <= memory2[ 3]; turn15 <= memory2[ 2]; 
					turn16 <= memory2[ 1]; turn17 <= memory2[ 0]; turn18 <= memory2[ 0]; 
				end
				2'd2: begin
					turn1 <= memory3[16]; turn2 <= memory3[15]; turn3 <= memory3[14]; 
					turn4 <= memory3[13]; turn5 <= memory3[12]; turn6 <= memory3[11]; 
					turn7 <= memory3[10]; turn8 <= memory3[ 9]; turn9 <= memory3[ 8]; 
					turn10 <= memory3[ 7]; turn11 <= memory3[ 6]; turn12 <= memory3[ 5]; 
					turn13 <= memory3[ 4]; turn14 <= memory3[ 3]; turn15 <= memory3[ 2]; 
					turn16 <= memory3[ 1]; turn17 <= memory3[ 0]; turn18 <= memory3[ 0]; 
				end
				2'd3: begin
					turn1 <= memory4[16]; turn2 <= memory4[15]; turn3 <= memory4[14]; 
					turn4 <= memory4[13]; turn5 <= memory4[12]; turn6 <= memory4[11]; 
					turn7 <= memory4[10]; turn8 <= memory4[ 9]; turn9 <= memory4[ 8]; 
					turn10 <= memory4[ 7]; turn11 <= memory4[ 6]; turn12 <= memory4[ 5]; 
					turn13 <= memory4[ 4]; turn14 <= memory4[ 3]; turn15 <= memory4[ 2]; 
					turn16 <= memory4[ 1]; turn17 <= memory4[ 0]; turn18 <= memory4[ 0]; 
				end
			endcase
        end else begin
            if(shift_enable) begin
                case(song)
                    2'd0: turn1 <= memory[cnt];
                    2'd1: turn1 <= memory2[cnt];
                    2'd2: turn1 <= memory3[cnt];
                    2'd3: turn1 <= memory4[cnt];                    
                endcase
				turn2 <= turn1; turn3 <= turn2; turn4 <= turn3; 
				turn5 <= turn4; turn6 <= turn5; turn7 <= turn6; 
				turn8 <= turn7; turn9 <= turn8; turn10 <= turn9; 
				turn11 <= turn10; turn12 <= turn11; turn13 <= turn12; 
				turn14 <= turn13; turn15 <= turn14; turn16 <= turn15; 
				turn17 <= turn16; turn18 <= turn17; 
            end
        end
    end
    // cnt for memory read address control
    always @(posedge clk or posedge reset) begin
        if(reset) begin
            cnt <= 17;
        end else begin 
            cnt <= cnt_next;
        end 
    end
    always@(*)begin
        if(load) begin
            cnt_next = 17;
        end else begin
            if(shift_enable) begin
                cnt_next = cnt + 1;
            end else begin
                cnt_next = cnt;
            end
        end
    end
    // ────────────────────────────────────────────────────────────────────────────────

    //
    // ─── JUDGE ROAD DISPLAY ─────────────────────────────────────────────────────────
    //

	assign is_road = (scan_in_turn12 | scan_in_turn23 | scan_in_turn34 | 
		scan_in_turn45 | scan_in_turn56 | scan_in_turn67 | scan_in_turn78 | 
		scan_in_turn89 | scan_in_turn910 | scan_in_turn1011 | scan_in_turn1112 | 
		scan_in_turn1213 | scan_in_turn1314 | scan_in_turn1415 | scan_in_turn1516 | 
		scan_in_turn1617 | scan_in_turn1718);

	assign scan_in_turn12 = 
    (
        turn1[10:0]==turn2[10:0] ? (current_block_x >= turn2[21:11] && current_block_x <= turn1[21:11])
        && current_block_y == turn1[10:0]
        : (current_block_y >= turn2[10:0] && current_block_y <= turn1[10:0])
        && current_block_x == turn1[21:11]
    );
	assign scan_in_turn23 = 
    (
        turn2[10:0]==turn3[10:0] ? (current_block_x >= turn3[21:11] && current_block_x <= turn2[21:11])
        && current_block_y == turn2[10:0]
        : (current_block_y >= turn3[10:0] && current_block_y <= turn2[10:0])
        && current_block_x == turn2[21:11]
    );
	assign scan_in_turn34 = 
    (
        turn3[10:0]==turn4[10:0] ? (current_block_x >= turn4[21:11] && current_block_x <= turn3[21:11])
        && current_block_y == turn3[10:0]
        : (current_block_y >= turn4[10:0] && current_block_y <= turn3[10:0])
        && current_block_x == turn3[21:11]
    );
	assign scan_in_turn45 = 
    (
        turn4[10:0]==turn5[10:0] ? (current_block_x >= turn5[21:11] && current_block_x <= turn4[21:11])
        && current_block_y == turn4[10:0]
        : (current_block_y >= turn5[10:0] && current_block_y <= turn4[10:0])
        && current_block_x == turn4[21:11]
    );
	assign scan_in_turn56 = 
    (
        turn5[10:0]==turn6[10:0] ? (current_block_x >= turn6[21:11] && current_block_x <= turn5[21:11])
        && current_block_y == turn5[10:0]
        : (current_block_y >= turn6[10:0] && current_block_y <= turn5[10:0])
        && current_block_x == turn5[21:11]
    );
	assign scan_in_turn67 = 
    (
        turn6[10:0]==turn7[10:0] ? (current_block_x >= turn7[21:11] && current_block_x <= turn6[21:11])
        && current_block_y == turn6[10:0]
        : (current_block_y >= turn7[10:0] && current_block_y <= turn6[10:0])
        && current_block_x == turn6[21:11]
    );
	assign scan_in_turn78 = 
    (
        turn7[10:0]==turn8[10:0] ? (current_block_x >= turn8[21:11] && current_block_x <= turn7[21:11])
        && current_block_y == turn7[10:0]
        : (current_block_y >= turn8[10:0] && current_block_y <= turn7[10:0])
        && current_block_x == turn7[21:11]
    );
	assign scan_in_turn89 = 
    (
        turn8[10:0]==turn9[10:0] ? (current_block_x >= turn9[21:11] && current_block_x <= turn8[21:11])
        && current_block_y == turn8[10:0]
        : (current_block_y >= turn9[10:0] && current_block_y <= turn8[10:0])
        && current_block_x == turn8[21:11]
    );
	assign scan_in_turn910 = 
    (
        turn9[10:0]==turn10[10:0] ? (current_block_x >= turn10[21:11] && current_block_x <= turn9[21:11])
        && current_block_y == turn9[10:0]
        : (current_block_y >= turn10[10:0] && current_block_y <= turn9[10:0])
        && current_block_x == turn9[21:11]
    );
	assign scan_in_turn1011 = 
    (
        turn10[10:0]==turn11[10:0] ? (current_block_x >= turn11[21:11] && current_block_x <= turn10[21:11])
        && current_block_y == turn10[10:0]
        : (current_block_y >= turn11[10:0] && current_block_y <= turn10[10:0])
        && current_block_x == turn10[21:11]
    );
	assign scan_in_turn1112 = 
    (
        turn11[10:0]==turn12[10:0] ? (current_block_x >= turn12[21:11] && current_block_x <= turn11[21:11])
        && current_block_y == turn11[10:0]
        : (current_block_y >= turn12[10:0] && current_block_y <= turn11[10:0])
        && current_block_x == turn11[21:11]
    );
	assign scan_in_turn1213 = 
    (
        turn12[10:0]==turn13[10:0] ? (current_block_x >= turn13[21:11] && current_block_x <= turn12[21:11])
        && current_block_y == turn12[10:0]
        : (current_block_y >= turn13[10:0] && current_block_y <= turn12[10:0])
        && current_block_x == turn12[21:11]
    );
	assign scan_in_turn1314 = 
    (
        turn13[10:0]==turn14[10:0] ? (current_block_x >= turn14[21:11] && current_block_x <= turn13[21:11])
        && current_block_y == turn13[10:0]
        : (current_block_y >= turn14[10:0] && current_block_y <= turn13[10:0])
        && current_block_x == turn13[21:11]
    );
	assign scan_in_turn1415 = 
    (
        turn14[10:0]==turn15[10:0] ? (current_block_x >= turn15[21:11] && current_block_x <= turn14[21:11])
        && current_block_y == turn14[10:0]
        : (current_block_y >= turn15[10:0] && current_block_y <= turn14[10:0])
        && current_block_x == turn14[21:11]
    );
	assign scan_in_turn1516 = 
    (
        turn15[10:0]==turn16[10:0] ? (current_block_x >= turn16[21:11] && current_block_x <= turn15[21:11])
        && current_block_y == turn15[10:0]
        : (current_block_y >= turn16[10:0] && current_block_y <= turn15[10:0])
        && current_block_x == turn15[21:11]
    );
	assign scan_in_turn1617 = 
    (
        turn16[10:0]==turn17[10:0] ? (current_block_x >= turn17[21:11] && current_block_x <= turn16[21:11])
        && current_block_y == turn16[10:0]
        : (current_block_y >= turn17[10:0] && current_block_y <= turn16[10:0])
        && current_block_x == turn16[21:11]
    );
	assign scan_in_turn1718 = 
    (
        turn17[10:0]==turn18[10:0] ? (current_block_x >= turn18[21:11] && current_block_x <= turn17[21:11])
        && current_block_y == turn17[10:0]
        : (current_block_y >= turn18[10:0] && current_block_y <= turn17[10:0])
        && current_block_x == turn17[21:11]
    );
    // ────────────────────────────────────────────────────────────────────────────────

    //
    // ─── JUDGE FAILED DISPLAY ───────────────────────────────────────────────────────
    //

    always@(posedge clk) begin
     fail = 
        ~(
            (dot1_in_turn12 | dot1_in_turn23 | dot1_in_turn34 | 
            dot1_in_turn45 | dot1_in_turn56 | dot1_in_turn67 | dot1_in_turn78 | 
            dot1_in_turn89 | dot1_in_turn910 | dot1_in_turn1011 | dot1_in_turn1112 | 
            dot1_in_turn1213 | dot1_in_turn1314 | dot1_in_turn1415 | dot1_in_turn1516 | 
            dot1_in_turn1617 | dot1_in_turn1718) | 
            (dot2_in_turn12 | dot2_in_turn23 | dot2_in_turn34 | 
            dot2_in_turn45 | dot2_in_turn56 | dot2_in_turn67 | dot2_in_turn78 | 
            dot2_in_turn89 | dot2_in_turn910 | dot2_in_turn1011 | dot2_in_turn1112 | 
            dot2_in_turn1213 | dot2_in_turn1314 | dot2_in_turn1415 | dot2_in_turn1516 | 
            dot2_in_turn1617 | dot2_in_turn1718) | 
            shift_enable 
        );
    end

    
    assign dot1_in_turn12 = (x1 >= turn2[21:11] && x1 <= turn1[21:11] && y1 >= turn2[10:0] && y1 <= turn1[10:0]);
    assign dot1_in_turn23 = (x1 >= turn3[21:11] && x1 <= turn2[21:11] && y1 >= turn3[10:0] && y1 <= turn2[10:0]);
    assign dot1_in_turn34 = (x1 >= turn4[21:11] && x1 <= turn3[21:11] && y1 >= turn4[10:0] && y1 <= turn3[10:0]);
    assign dot1_in_turn45 = (x1 >= turn5[21:11] && x1 <= turn4[21:11] && y1 >= turn5[10:0] && y1 <= turn4[10:0]);
    assign dot1_in_turn56 = (x1 >= turn6[21:11] && x1 <= turn5[21:11] && y1 >= turn6[10:0] && y1 <= turn5[10:0]);
    assign dot1_in_turn67 = (x1 >= turn7[21:11] && x1 <= turn6[21:11] && y1 >= turn7[10:0] && y1 <= turn6[10:0]);
    assign dot1_in_turn78 = (x1 >= turn8[21:11] && x1 <= turn7[21:11] && y1 >= turn8[10:0] && y1 <= turn7[10:0]);
    assign dot1_in_turn89 = (x1 >= turn9[21:11] && x1 <= turn8[21:11] && y1 >= turn9[10:0] && y1 <= turn8[10:0]);
    assign dot1_in_turn910 = (x1 >= turn10[21:11] && x1 <= turn9[21:11] && y1 >= turn10[10:0] && y1 <= turn9[10:0]);
    assign dot1_in_turn1011 = (x1 >= turn11[21:11] && x1 <= turn10[21:11] && y1 >= turn11[10:0] && y1 <= turn10[10:0]);
    assign dot1_in_turn1112 = (x1 >= turn12[21:11] && x1 <= turn11[21:11] && y1 >= turn12[10:0] && y1 <= turn11[10:0]);
    assign dot1_in_turn1213 = (x1 >= turn13[21:11] && x1 <= turn12[21:11] && y1 >= turn13[10:0] && y1 <= turn12[10:0]);
    assign dot1_in_turn1314 = (x1 >= turn14[21:11] && x1 <= turn13[21:11] && y1 >= turn14[10:0] && y1 <= turn13[10:0]);
    assign dot1_in_turn1415 = (x1 >= turn15[21:11] && x1 <= turn14[21:11] && y1 >= turn15[10:0] && y1 <= turn14[10:0]);
    assign dot1_in_turn1516 = (x1 >= turn16[21:11] && x1 <= turn15[21:11] && y1 >= turn16[10:0] && y1 <= turn15[10:0]);
    assign dot1_in_turn1617 = (x1 >= turn17[21:11] && x1 <= turn16[21:11] && y1 >= turn17[10:0] && y1 <= turn16[10:0]);
    assign dot1_in_turn1718 = (x1 >= turn18[21:11] && x1 <= turn17[21:11] && y1 >= turn18[10:0] && y1 <= turn17[10:0]);
    assign dot2_in_turn12 = (x2 >= turn2[21:11] && x2 <= turn1[21:11] && y2 >= turn2[10:0] && y2 <= turn1[10:0]);
    assign dot2_in_turn23 = (x2 >= turn3[21:11] && x2 <= turn2[21:11] && y2 >= turn3[10:0] && y2 <= turn2[10:0]);
    assign dot2_in_turn34 = (x2 >= turn4[21:11] && x2 <= turn3[21:11] && y2 >= turn4[10:0] && y2 <= turn3[10:0]);
    assign dot2_in_turn45 = (x2 >= turn5[21:11] && x2 <= turn4[21:11] && y2 >= turn5[10:0] && y2 <= turn4[10:0]);
    assign dot2_in_turn56 = (x2 >= turn6[21:11] && x2 <= turn5[21:11] && y2 >= turn6[10:0] && y2 <= turn5[10:0]);
    assign dot2_in_turn67 = (x2 >= turn7[21:11] && x2 <= turn6[21:11] && y2 >= turn7[10:0] && y2 <= turn6[10:0]);
    assign dot2_in_turn78 = (x2 >= turn8[21:11] && x2 <= turn7[21:11] && y2 >= turn8[10:0] && y2 <= turn7[10:0]);
    assign dot2_in_turn89 = (x2 >= turn9[21:11] && x2 <= turn8[21:11] && y2 >= turn9[10:0] && y2 <= turn8[10:0]);
    assign dot2_in_turn910 = (x2 >= turn10[21:11] && x2 <= turn9[21:11] && y2 >= turn10[10:0] && y2 <= turn9[10:0]);
    assign dot2_in_turn1011 = (x2 >= turn11[21:11] && x2 <= turn10[21:11] && y2 >= turn11[10:0] && y2 <= turn10[10:0]);
    assign dot2_in_turn1112 = (x2 >= turn12[21:11] && x2 <= turn11[21:11] && y2 >= turn12[10:0] && y2 <= turn11[10:0]);
    assign dot2_in_turn1213 = (x2 >= turn13[21:11] && x2 <= turn12[21:11] && y2 >= turn13[10:0] && y2 <= turn12[10:0]);
    assign dot2_in_turn1314 = (x2 >= turn14[21:11] && x2 <= turn13[21:11] && y2 >= turn14[10:0] && y2 <= turn13[10:0]);
    assign dot2_in_turn1415 = (x2 >= turn15[21:11] && x2 <= turn14[21:11] && y2 >= turn15[10:0] && y2 <= turn14[10:0]);
    assign dot2_in_turn1516 = (x2 >= turn16[21:11] && x2 <= turn15[21:11] && y2 >= turn16[10:0] && y2 <= turn15[10:0]);
    assign dot2_in_turn1617 = (x2 >= turn17[21:11] && x2 <= turn16[21:11] && y2 >= turn17[10:0] && y2 <= turn16[10:0]);
    assign dot2_in_turn1718 = (x2 >= turn18[21:11] && x2 <= turn17[21:11] && y2 >= turn18[10:0] && y2 <= turn17[10:0]);
    // ────────────────────────────────────────────────────────────────────────────────

    //
    // ─── COORDINATES ────────────────────────────────────────────────────────────────
    //
    //                   (       x,       y)
    assign memory[  0] = {11'd  10,11'd   7};
    assign memory[  1] = {11'd  14,11'd   7};
    assign memory[  2] = {11'd  14,11'd  15};
    assign memory[  3] = {11'd  22,11'd  15};
    assign memory[  4] = {11'd  22,11'd  23};
    assign memory[  5] = {11'd  30,11'd  23};
    assign memory[  6] = {11'd  30,11'd  31};
    assign memory[  7] = {11'd  34,11'd  31};
    assign memory[  8] = {11'd  34,11'd  34};
    assign memory[  9] = {11'd  37,11'd  34};
    assign memory[ 10] = {11'd  37,11'd  36};
    assign memory[ 11] = {11'd  41,11'd  36};
    assign memory[ 12] = {11'd  41,11'd  40};
    assign memory[ 13] = {11'd  45,11'd  40};
    assign memory[ 14] = {11'd  45,11'd  44};
    assign memory[ 15] = {11'd  49,11'd  44};
    assign memory[ 16] = {11'd  49,11'd  48};
    assign memory[ 17] = {11'd  51,11'd  48};
    assign memory[ 18] = {11'd  51,11'd  50};
    assign memory[ 19] = {11'd  53,11'd  50};
    assign memory[ 20] = {11'd  53,11'd  52};
    assign memory[ 21] = {11'd  57,11'd  52};
    assign memory[ 22] = {11'd  57,11'd  56};
    assign memory[ 23] = {11'd  61,11'd  56};
    assign memory[ 24] = {11'd  61,11'd  60};
    assign memory[ 25] = {11'd  63,11'd  60};
    assign memory[ 26] = {11'd  63,11'd  62};
    assign memory[ 27] = {11'd  65,11'd  62};
    assign memory[ 28] = {11'd  65,11'd  64};
    assign memory[ 29] = {11'd  69,11'd  64};
    assign memory[ 30] = {11'd  69,11'd  68};
    assign memory[ 31] = {11'd  71,11'd  68};
    assign memory[ 32] = {11'd  71,11'd  70};
    assign memory[ 33] = {11'd  73,11'd  70};
    assign memory[ 34] = {11'd  73,11'd  72};
    assign memory[ 35] = {11'd  77,11'd  72};
    assign memory[ 36] = {11'd  77,11'd  76};
    assign memory[ 37] = {11'd  83,11'd  76};
    assign memory[ 38] = {11'd  83,11'd  78};
    assign memory[ 39] = {11'd  87,11'd  78};
    assign memory[ 40] = {11'd  87,11'd  82};
    assign memory[ 41] = {11'd  89,11'd  82};
    assign memory[ 42] = {11'd  89,11'd  84};
    assign memory[ 43] = {11'd  91,11'd  84};
    assign memory[ 44] = {11'd  91,11'd  86};
    assign memory[ 45] = {11'd  93,11'd  86};
    assign memory[ 46] = {11'd  93,11'd  88};
    assign memory[ 47] = {11'd  95,11'd  88};
    assign memory[ 48] = {11'd  95,11'd  90};
    assign memory[ 49] = {11'd  97,11'd  90};
    assign memory[ 50] = {11'd  97,11'd  92};
    assign memory[ 51] = {11'd  99,11'd  92};
    assign memory[ 52] = {11'd  99,11'd  94};
    assign memory[ 53] = {11'd 111,11'd  94};
    assign memory[ 54] = {11'd 111,11'd  98};
    assign memory[ 55] = {11'd 115,11'd  98};
    assign memory[ 56] = {11'd 115,11'd 102};
    assign memory[ 57] = {11'd 119,11'd 102};
    assign memory[ 58] = {11'd 119,11'd 106};
    assign memory[ 59] = {11'd 121,11'd 106};
    assign memory[ 60] = {11'd 121,11'd 108};
    assign memory[ 61] = {11'd 123,11'd 108};
    assign memory[ 62] = {11'd 123,11'd 110};
    assign memory[ 63] = {11'd 127,11'd 110};
    assign memory[ 64] = {11'd 127,11'd 114};
    assign memory[ 65] = {11'd 131,11'd 114};
    assign memory[ 66] = {11'd 131,11'd 118};
    assign memory[ 67] = {11'd 135,11'd 118};
    assign memory[ 68] = {11'd 135,11'd 122};
    assign memory[ 69] = {11'd 137,11'd 122};
    assign memory[ 70] = {11'd 137,11'd 124};
    assign memory[ 71] = {11'd 139,11'd 124};
    assign memory[ 72] = {11'd 139,11'd 126};
    assign memory[ 73] = {11'd 143,11'd 126};
    assign memory[ 74] = {11'd 143,11'd 128};
    assign memory[ 75] = {11'd 145,11'd 128};
    assign memory[ 76] = {11'd 145,11'd 132};
    assign memory[ 77] = {11'd 149,11'd 132};
    assign memory[ 78] = {11'd 149,11'd 136};
    assign memory[ 79] = {11'd 153,11'd 136};
    assign memory[ 80] = {11'd 153,11'd 138};
    assign memory[ 81] = {11'd 155,11'd 138};
    assign memory[ 82] = {11'd 155,11'd 140};
    assign memory[ 83] = {11'd 157,11'd 140};
    assign memory[ 84] = {11'd 157,11'd 144};
    assign memory[ 85] = {11'd 161,11'd 144};
    assign memory[ 86] = {11'd 161,11'd 148};
    assign memory[ 87] = {11'd 165,11'd 148};
    assign memory[ 88] = {11'd 165,11'd 150};
    assign memory[ 89] = {11'd 167,11'd 150};
    assign memory[ 90] = {11'd 167,11'd 152};
    assign memory[ 91] = {11'd 169,11'd 152};
    assign memory[ 92] = {11'd 169,11'd 164};
    assign memory[ 93] = {11'd 173,11'd 164};
    assign memory[ 94] = {11'd 173,11'd 168};
    assign memory[ 95] = {11'd 175,11'd 168};
    assign memory[ 96] = {11'd 175,11'd 170};
    assign memory[ 97] = {11'd 179,11'd 170};
    assign memory[ 98] = {11'd 179,11'd 172};
    assign memory[ 99] = {11'd 181,11'd 172};
    assign memory[100] = {11'd 181,11'd 174};
    assign memory[101] = {11'd 183,11'd 174};
    assign memory[102] = {11'd 183,11'd 176};
    assign memory[103] = {11'd 185,11'd 176};
    assign memory[104] = {11'd 185,11'd 180};
    assign memory[105] = {11'd 189,11'd 180};
    assign memory[106] = {11'd 189,11'd 184};
    assign memory[107] = {11'd 191,11'd 184};
    assign memory[108] = {11'd 191,11'd 186};
    assign memory[109] = {11'd 195,11'd 186};
    assign memory[110] = {11'd 195,11'd 188};
    assign memory[111] = {11'd 197,11'd 188};
    assign memory[112] = {11'd 197,11'd 190};
    assign memory[113] = {11'd 199,11'd 190};
    assign memory[114] = {11'd 199,11'd 192};
    assign memory[115] = {11'd 201,11'd 192};
    assign memory[116] = {11'd 201,11'd 196};
    assign memory[117] = {11'd 203,11'd 196};
    assign memory[118] = {11'd 203,11'd 198};
    assign memory[119] = {11'd 207,11'd 198};
    assign memory[120] = {11'd 207,11'd 200};
    assign memory[121] = {11'd 209,11'd 200};
    assign memory[122] = {11'd 209,11'd 202};
    assign memory[123] = {11'd 211,11'd 202};
    assign memory[124] = {11'd 211,11'd 204};
    assign memory[125] = {11'd 213,11'd 204};
    assign memory[126] = {11'd 213,11'd 206};
    assign memory[127] = {11'd 215,11'd 206};
    assign memory[128] = {11'd 215,11'd 208};
    assign memory[129] = {11'd 217,11'd 208};
    assign memory[130] = {11'd 217,11'd 212};
    assign memory[131] = {11'd 221,11'd 212};
    assign memory[132] = {11'd 221,11'd 216};
    assign memory[133] = {11'd 223,11'd 216};
    assign memory[134] = {11'd 223,11'd 218};
    assign memory[135] = {11'd 225,11'd 218};
    assign memory[136] = {11'd 225,11'd 220};
    assign memory[137] = {11'd 227,11'd 220};
    assign memory[138] = {11'd 227,11'd 222};
    assign memory[139] = {11'd 239,11'd 222};
    assign memory[140] = {11'd 239,11'd 226};
    assign memory[141] = {11'd 247,11'd 226};
    assign memory[142] = {11'd 247,11'd 234};
    assign memory[143] = {11'd 255,11'd 234};
    assign memory[144] = {11'd 255,11'd 242};
    assign memory[145] = {11'd 267,11'd 242};
    assign memory[146] = {11'd 267,11'd 246};
    assign memory[147] = {11'd 275,11'd 246};
    assign memory[148] = {11'd 275,11'd 250};
    assign memory[149] = {11'd 279,11'd 250};
    assign memory[150] = {11'd 279,11'd 258};
    assign memory[151] = {11'd 287,11'd 258};
    assign memory[152] = {11'd 287,11'd 266};
    assign memory[153] = {11'd 295,11'd 266};
    assign memory[154] = {11'd 295,11'd 278};
    assign memory[155] = {11'd 299,11'd 278};
    assign memory[156] = {11'd 299,11'd 282};
    assign memory[157] = {11'd 303,11'd 282};
    assign memory[158] = {11'd 303,11'd 286};
    assign memory[159] = {11'd 307,11'd 286};
    assign memory[160] = {11'd 307,11'd 294};
    assign memory[161] = {11'd 315,11'd 294};
    assign memory[162] = {11'd 315,11'd 302};
    assign memory[163] = {11'd 323,11'd 302};
    assign memory[164] = {11'd 323,11'd 314};
    assign memory[165] = {11'd 327,11'd 314};
    assign memory[166] = {11'd 327,11'd 322};
    assign memory[167] = {11'd 331,11'd 322};
    assign memory[168] = {11'd 331,11'd 326};
    assign memory[169] = {11'd 339,11'd 326};
    assign memory[170] = {11'd 339,11'd 334};
    assign memory[171] = {11'd 347,11'd 334};
    assign memory[172] = {11'd 347,11'd 342};
    assign memory[173] = {11'd 359,11'd 342};
    assign memory[174] = {11'd 359,11'd 346};
    assign memory[175] = {11'd 363,11'd 346};
    assign memory[176] = {11'd 363,11'd 350};
    assign memory[177] = {11'd 367,11'd 350};
    assign memory[178] = {11'd 367,11'd 358};
    assign memory[179] = {11'd 375,11'd 358};
    assign memory[180] = {11'd 375,11'd 366};
    assign memory[181] = {11'd 383,11'd 366};
    assign memory[182] = {11'd 383,11'd 374};
    assign memory[183] = {11'd 391,11'd 374};
    assign memory[184] = {11'd 391,11'd 378};
    assign memory[185] = {11'd 394,11'd 378};
    assign memory[186] = {11'd 394,11'd 381};
    assign memory[187] = {11'd 396,11'd 381};
    assign memory[188] = {11'd 396,11'd 389};
    assign memory[189] = {11'd 400,11'd 389};
    assign memory[190] = {11'd 400,11'd 391};
    assign memory[191] = {11'd 402,11'd 391};
    assign memory[192] = {11'd 402,11'd 395};
    assign memory[193] = {11'd 404,11'd 395};
    assign memory[194] = {11'd 404,11'd 397};
    assign memory[195] = {11'd 406,11'd 397};
    assign memory[196] = {11'd 406,11'd 399};
    assign memory[197] = {11'd 408,11'd 399};
    assign memory[198] = {11'd 408,11'd 401};
    assign memory[199] = {11'd 412,11'd 401};
    assign memory[200] = {11'd 412,11'd 403};
    assign memory[201] = {11'd 414,11'd 403};
    assign memory[202] = {11'd 414,11'd 407};
    assign memory[203] = {11'd 416,11'd 407};
    assign memory[204] = {11'd 416,11'd 409};
    assign memory[205] = {11'd 418,11'd 409};
    assign memory[206] = {11'd 418,11'd 411};
    assign memory[207] = {11'd 420,11'd 411};
    assign memory[208] = {11'd 420,11'd 413};
    assign memory[209] = {11'd 424,11'd 413};
    assign memory[210] = {11'd 424,11'd 415};
    assign memory[211] = {11'd 426,11'd 415};
    assign memory[212] = {11'd 426,11'd 417};
    assign memory[213] = {11'd 428,11'd 417};
    assign memory[214] = {11'd 428,11'd 419};
    assign memory[215] = {11'd 430,11'd 419};
    assign memory[216] = {11'd 430,11'd 421};
    assign memory[217] = {11'd 432,11'd 421};
    assign memory[218] = {11'd 432,11'd 423};
    assign memory[219] = {11'd 434,11'd 423};
    assign memory[220] = {11'd 434,11'd 429};
    assign memory[221] = {11'd 436,11'd 429};
    assign memory[222] = {11'd 436,11'd 433};
    assign memory[223] = {11'd 440,11'd 433};
    assign memory[224] = {11'd 440,11'd 435};
    assign memory[225] = {11'd 442,11'd 435};
    assign memory[226] = {11'd 442,11'd 437};
    assign memory[227] = {11'd 444,11'd 437};
    assign memory[228] = {11'd 444,11'd 439};
    assign memory[229] = {11'd 446,11'd 439};
    assign memory[230] = {11'd 446,11'd 441};
    assign memory[231] = {11'd 448,11'd 441};
    assign memory[232] = {11'd 448,11'd 443};
    assign memory[233] = {11'd 450,11'd 443};
    assign memory[234] = {11'd 450,11'd 445};
    assign memory[235] = {11'd 452,11'd 445};
    assign memory[236] = {11'd 452,11'd 457};
    assign memory[237] = {11'd 456,11'd 457};
    assign memory[238] = {11'd 456,11'd 461};
    assign memory[239] = {11'd 458,11'd 461};
    assign memory[240] = {11'd 458,11'd 463};
    assign memory[241] = {11'd 462,11'd 463};
    assign memory[242] = {11'd 462,11'd 465};
    assign memory[243] = {11'd 464,11'd 465};
    assign memory[244] = {11'd 464,11'd 467};
    assign memory[245] = {11'd 466,11'd 467};
    assign memory[246] = {11'd 466,11'd 469};
    assign memory[247] = {11'd 468,11'd 469};
    assign memory[248] = {11'd 468,11'd 473};
    assign memory[249] = {11'd 472,11'd 473};
    assign memory[250] = {11'd 472,11'd 477};
    assign memory[251] = {11'd 474,11'd 477};
    assign memory[252] = {11'd 474,11'd 479};
    assign memory[253] = {11'd 478,11'd 479};
    assign memory[254] = {11'd 478,11'd 481};
    assign memory[255] = {11'd 480,11'd 481};
    assign memory[256] = {11'd 480,11'd 483};
    assign memory[257] = {11'd 482,11'd 483};
    assign memory[258] = {11'd 482,11'd 485};
    assign memory[259] = {11'd 484,11'd 485};
    assign memory[260] = {11'd 484,11'd 489};
    assign memory[261] = {11'd 486,11'd 489};
    assign memory[262] = {11'd 486,11'd 491};
    assign memory[263] = {11'd 490,11'd 491};
    assign memory[264] = {11'd 490,11'd 493};
    assign memory[265] = {11'd 492,11'd 493};
    assign memory[266] = {11'd 492,11'd 495};
    assign memory[267] = {11'd 494,11'd 495};
    assign memory[268] = {11'd 494,11'd 497};
    assign memory[269] = {11'd 496,11'd 497};
    assign memory[270] = {11'd 496,11'd 499};
    assign memory[271] = {11'd 498,11'd 499};
    assign memory[272] = {11'd 498,11'd 501};
    assign memory[273] = {11'd 500,11'd 501};
    assign memory[274] = {11'd 500,11'd 505};
    assign memory[275] = {11'd 504,11'd 505};
    assign memory[276] = {11'd 504,11'd 509};
    assign memory[277] = {11'd 506,11'd 509};
    assign memory[278] = {11'd 506,11'd 511};
    assign memory[279] = {11'd 508,11'd 511};
    assign memory[280] = {11'd 508,11'd 513};
    assign memory[281] = {11'd 510,11'd 513};
    assign memory[282] = {11'd 510,11'd 515};
    assign memory[283] = {11'd 522,11'd 515};
    assign memory[284] = {11'd 522,11'd 517};
    assign memory[285] = {11'd 524,11'd 517};
    assign memory[286] = {11'd 524,11'd 521};
    assign memory[287] = {11'd 526,11'd 521};
    assign memory[288] = {11'd 526,11'd 523};
    assign memory[289] = {11'd 530,11'd 523};
    assign memory[290] = {11'd 530,11'd 525};
    assign memory[291] = {11'd 532,11'd 525};
    assign memory[292] = {11'd 532,11'd 527};
    assign memory[293] = {11'd 534,11'd 527};
    assign memory[294] = {11'd 534,11'd 529};
    assign memory[295] = {11'd 536,11'd 529};
    assign memory[296] = {11'd 536,11'd 533};
    assign memory[297] = {11'd 540,11'd 533};
    assign memory[298] = {11'd 540,11'd 537};
    assign memory[299] = {11'd 542,11'd 537};
    assign memory[300] = {11'd 542,11'd 539};
    assign memory[301] = {11'd 544,11'd 539};
    assign memory[302] = {11'd 544,11'd 541};
    assign memory[303] = {11'd 546,11'd 541};
    assign memory[304] = {11'd 546,11'd 543};
    assign memory[305] = {11'd 548,11'd 543};
    assign memory[306] = {11'd 548,11'd 545};
    assign memory[307] = {11'd 550,11'd 545};
    assign memory[308] = {11'd 550,11'd 547};
    assign memory[309] = {11'd 554,11'd 547};
    assign memory[310] = {11'd 554,11'd 549};
    assign memory[311] = {11'd 556,11'd 549};
    assign memory[312] = {11'd 556,11'd 553};
    assign memory[313] = {11'd 558,11'd 553};
    assign memory[314] = {11'd 558,11'd 555};
    assign memory[315] = {11'd 560,11'd 555};
    assign memory[316] = {11'd 560,11'd 557};
    assign memory[317] = {11'd 562,11'd 557};
    assign memory[318] = {11'd 562,11'd 559};
    assign memory[319] = {11'd 564,11'd 559};
    assign memory[320] = {11'd 564,11'd 561};
    assign memory[321] = {11'd 566,11'd 561};
    assign memory[322] = {11'd 566,11'd 563};
    assign memory[323] = {11'd 570,11'd 563};
    assign memory[324] = {11'd 570,11'd 567};
    assign memory[325] = {11'd 574,11'd 567};
    assign memory[326] = {11'd 574,11'd 569};
    assign memory[327] = {11'd 576,11'd 569};
    assign memory[328] = {11'd 576,11'd 571};
    assign memory[329] = {11'd 578,11'd 571};
    assign memory[330] = {11'd 578,11'd 573};
    assign memory[331] = {11'd 580,11'd 573};
    assign memory[332] = {11'd 580,11'd 585};
    assign memory[333] = {11'd 582,11'd 585};
    assign memory[334] = {11'd 582,11'd 587};
    assign memory[335] = {11'd 586,11'd 587};
    assign memory[336] = {11'd 586,11'd 589};
    assign memory[337] = {11'd 588,11'd 589};
    assign memory[338] = {11'd 588,11'd 593};
    assign memory[339] = {11'd 590,11'd 593};
    assign memory[340] = {11'd 590,11'd 595};
    assign memory[341] = {11'd 592,11'd 595};
    assign memory[342] = {11'd 592,11'd 597};
    assign memory[343] = {11'd 594,11'd 597};
    assign memory[344] = {11'd 594,11'd 599};
    assign memory[345] = {11'd 598,11'd 599};
    assign memory[346] = {11'd 598,11'd 601};
    assign memory[347] = {11'd 600,11'd 601};
    assign memory[348] = {11'd 600,11'd 605};
    assign memory[349] = {11'd 602,11'd 605};
    assign memory[350] = {11'd 602,11'd 607};
    assign memory[351] = {11'd 604,11'd 607};
    assign memory[352] = {11'd 604,11'd 609};
    assign memory[353] = {11'd 606,11'd 609};
    assign memory[354] = {11'd 606,11'd 611};
    assign memory[355] = {11'd 608,11'd 611};
    assign memory[356] = {11'd 608,11'd 613};
    assign memory[357] = {11'd 610,11'd 613};
    assign memory[358] = {11'd 610,11'd 615};
    assign memory[359] = {11'd 614,11'd 615};
    assign memory[360] = {11'd 614,11'd 617};
    assign memory[361] = {11'd 616,11'd 617};
    assign memory[362] = {11'd 616,11'd 621};
    assign memory[363] = {11'd 618,11'd 621};
    assign memory[364] = {11'd 618,11'd 623};
    assign memory[365] = {11'd 620,11'd 623};
    assign memory[366] = {11'd 620,11'd 625};
    assign memory[367] = {11'd 622,11'd 625};
    assign memory[368] = {11'd 622,11'd 627};
    assign memory[369] = {11'd 624,11'd 627};
    assign memory[370] = {11'd 624,11'd 629};
    assign memory[371] = {11'd 626,11'd 629};
    assign memory[372] = {11'd 626,11'd 631};
    assign memory[373] = {11'd 630,11'd 631};
    assign memory[374] = {11'd 630,11'd 633};
    assign memory[375] = {11'd 632,11'd 633};
    assign memory[376] = {11'd 632,11'd 637};
    assign memory[377] = {11'd 634,11'd 637};
    assign memory[378] = {11'd 634,11'd 639};
    assign memory[379] = {11'd 636,11'd 639};
    assign memory[380] = {11'd 636,11'd 641};
    assign memory[381] = {11'd 638,11'd 641};
    assign memory[382] = {11'd 638,11'd 643};
    assign memory[383] = {11'd 650,11'd 643};
    assign memory[384] = {11'd 650,11'd 645};
    assign memory[385] = {11'd 652,11'd 645};
    assign memory[386] = {11'd 652,11'd 649};
    assign memory[387] = {11'd 654,11'd 649};
    assign memory[388] = {11'd 654,11'd 651};
    assign memory[389] = {11'd 658,11'd 651};
    assign memory[390] = {11'd 658,11'd 653};
    assign memory[391] = {11'd 660,11'd 653};
    assign memory[392] = {11'd 660,11'd 655};
    assign memory[393] = {11'd 662,11'd 655};
    assign memory[394] = {11'd 662,11'd 657};
    assign memory[395] = {11'd 664,11'd 657};
    assign memory[396] = {11'd 664,11'd 661};
    assign memory[397] = {11'd 666,11'd 661};
    assign memory[398] = {11'd 666,11'd 663};
    assign memory[399] = {11'd 670,11'd 663};
    assign memory[400] = {11'd 670,11'd 665};
    assign memory[401] = {11'd 672,11'd 665};
    assign memory[402] = {11'd 672,11'd 667};
    assign memory[403] = {11'd 674,11'd 667};
    assign memory[404] = {11'd 674,11'd 669};
    assign memory[405] = {11'd 676,11'd 669};
    assign memory[406] = {11'd 676,11'd 671};
    assign memory[407] = {11'd 678,11'd 671};
    assign memory[408] = {11'd 678,11'd 673};
    assign memory[409] = {11'd 680,11'd 673};
    assign memory[410] = {11'd 680,11'd 677};
    assign memory[411] = {11'd 682,11'd 677};
    assign memory[412] = {11'd 682,11'd 679};
    assign memory[413] = {11'd 686,11'd 679};
    assign memory[414] = {11'd 686,11'd 681};
    assign memory[415] = {11'd 688,11'd 681};
    assign memory[416] = {11'd 688,11'd 683};
    assign memory[417] = {11'd 690,11'd 683};
    assign memory[418] = {11'd 690,11'd 685};
    assign memory[419] = {11'd 692,11'd 685};
    assign memory[420] = {11'd 692,11'd 687};
    assign memory[421] = {11'd 694,11'd 687};
    assign memory[422] = {11'd 694,11'd 689};
    assign memory[423] = {11'd 696,11'd 689};
    assign memory[424] = {11'd 696,11'd 693};
    assign memory[425] = {11'd 698,11'd 693};
    assign memory[426] = {11'd 698,11'd 695};
    assign memory[427] = {11'd 702,11'd 695};
    assign memory[428] = {11'd 702,11'd 697};
    assign memory[429] = {11'd 704,11'd 697};
    assign memory[430] = {11'd 704,11'd 699};
    assign memory[431] = {11'd 706,11'd 699};
    assign memory[432] = {11'd 706,11'd 701};
    assign memory[433] = {11'd 708,11'd 701};
    assign memory[434] = {11'd 708,11'd 713};
    assign memory[435] = {11'd 710,11'd 713};
    assign memory[436] = {11'd 710,11'd 715};
    assign memory[437] = {11'd 716,11'd 715};
    assign memory[438] = {11'd 716,11'd 717};
    assign memory[439] = {11'd 722,11'd 717};
    assign memory[440] = {11'd 722,11'd 719};
    assign memory[441] = {11'd 728,11'd 719};
    assign memory[442] = {11'd 728,11'd 721};
    assign memory[443] = {11'd 732,11'd 721};
    assign memory[444] = {11'd 732,11'd 725};
    assign memory[445] = {11'd 738,11'd 725};
    assign memory[446] = {11'd 738,11'd 727};
    assign memory[447] = {11'd 742,11'd 727};
    assign memory[448] = {11'd 742,11'd 731};
    assign memory[449] = {11'd 745,11'd 731};
    assign memory[450] = {11'd 745,11'd 734};
    assign memory[451] = {11'd 747,11'd 734};
    assign memory[452] = {11'd 747,11'd 742};
    assign memory[453] = {11'd 747,11'd 762};

    assign memory2[  0] = {11'd  10,11'd   7};
    assign memory2[  1] = {11'd  14,11'd   7};
    assign memory2[  2] = {11'd  14,11'd  11};
    assign memory2[  3] = {11'd  18,11'd  11};
    assign memory2[  4] = {11'd  18,11'd  15};
    assign memory2[  5] = {11'd  22,11'd  15};
    assign memory2[  6] = {11'd  22,11'd  19};
    assign memory2[  7] = {11'd  26,11'd  19};
    assign memory2[  8] = {11'd  26,11'd  23};
    assign memory2[  9] = {11'd  30,11'd  23};
    assign memory2[ 10] = {11'd  30,11'd  27};
    assign memory2[ 11] = {11'd  34,11'd  27};
    assign memory2[ 12] = {11'd  34,11'd  31};
    assign memory2[ 13] = {11'd  38,11'd  31};
    assign memory2[ 14] = {11'd  38,11'd  35};
    assign memory2[ 15] = {11'd  42,11'd  35};
    assign memory2[ 16] = {11'd  42,11'd  39};
    assign memory2[ 17] = {11'd  46,11'd  39};
    assign memory2[ 18] = {11'd  46,11'd  43};
    assign memory2[ 19] = {11'd  50,11'd  43};
    assign memory2[ 20] = {11'd  50,11'd  47};
    assign memory2[ 21] = {11'd  54,11'd  47};
    assign memory2[ 22] = {11'd  54,11'd  51};
    assign memory2[ 23] = {11'd  58,11'd  51};
    assign memory2[ 24] = {11'd  58,11'd  55};
    assign memory2[ 25] = {11'd  62,11'd  55};
    assign memory2[ 26] = {11'd  62,11'd  59};
    assign memory2[ 27] = {11'd  66,11'd  59};
    assign memory2[ 28] = {11'd  66,11'd  63};
    assign memory2[ 29] = {11'd  70,11'd  63};
    assign memory2[ 30] = {11'd  70,11'd  67};
    assign memory2[ 31] = {11'd  74,11'd  67};
    assign memory2[ 32] = {11'd  74,11'd  71};
    assign memory2[ 33] = {11'd  78,11'd  71};
    assign memory2[ 34] = {11'd  78,11'd  73};
    assign memory2[ 35] = {11'd  80,11'd  73};
    assign memory2[ 36] = {11'd  80,11'd  77};
    assign memory2[ 37] = {11'd  82,11'd  77};
    assign memory2[ 38] = {11'd  82,11'd  79};
    assign memory2[ 39] = {11'd  86,11'd  79};
    assign memory2[ 40] = {11'd  86,11'd  81};
    assign memory2[ 41] = {11'd  88,11'd  81};
    assign memory2[ 42] = {11'd  88,11'd  85};
    assign memory2[ 43] = {11'd  90,11'd  85};
    assign memory2[ 44] = {11'd  90,11'd  86};
    assign memory2[ 45] = {11'd  91,11'd  86};
    assign memory2[ 46] = {11'd  91,11'd  90};
    assign memory2[ 47] = {11'd  93,11'd  90};
    assign memory2[ 48] = {11'd  93,11'd  92};
    assign memory2[ 49] = {11'd  97,11'd  92};
    assign memory2[ 50] = {11'd  97,11'd  94};
    assign memory2[ 51] = {11'd  99,11'd  94};
    assign memory2[ 52] = {11'd  99,11'd  98};
    assign memory2[ 53] = {11'd 101,11'd  98};
    assign memory2[ 54] = {11'd 101,11'd 100};
    assign memory2[ 55] = {11'd 105,11'd 100};
    assign memory2[ 56] = {11'd 105,11'd 102};
    assign memory2[ 57] = {11'd 107,11'd 102};
    assign memory2[ 58] = {11'd 107,11'd 106};
    assign memory2[ 59] = {11'd 109,11'd 106};
    assign memory2[ 60] = {11'd 109,11'd 108};
    assign memory2[ 61] = {11'd 113,11'd 108};
    assign memory2[ 62] = {11'd 113,11'd 110};
    assign memory2[ 63] = {11'd 115,11'd 110};
    assign memory2[ 64] = {11'd 115,11'd 114};
    assign memory2[ 65] = {11'd 117,11'd 114};
    assign memory2[ 66] = {11'd 117,11'd 116};
    assign memory2[ 67] = {11'd 121,11'd 116};
    assign memory2[ 68] = {11'd 121,11'd 118};
    assign memory2[ 69] = {11'd 122,11'd 118};
    assign memory2[ 70] = {11'd 122,11'd 119};
    assign memory2[ 71] = {11'd 126,11'd 119};
    assign memory2[ 72] = {11'd 126,11'd 121};
    assign memory2[ 73] = {11'd 128,11'd 121};
    assign memory2[ 74] = {11'd 128,11'd 125};
    assign memory2[ 75] = {11'd 130,11'd 125};
    assign memory2[ 76] = {11'd 130,11'd 127};
    assign memory2[ 77] = {11'd 134,11'd 127};
    assign memory2[ 78] = {11'd 134,11'd 129};
    assign memory2[ 79] = {11'd 136,11'd 129};
    assign memory2[ 80] = {11'd 136,11'd 131};
    assign memory2[ 81] = {11'd 137,11'd 131};
    assign memory2[ 82] = {11'd 137,11'd 132};
    assign memory2[ 83] = {11'd 139,11'd 132};
    assign memory2[ 84] = {11'd 139,11'd 133};
    assign memory2[ 85] = {11'd 140,11'd 133};
    assign memory2[ 86] = {11'd 140,11'd 137};
    assign memory2[ 87] = {11'd 144,11'd 137};
    assign memory2[ 88] = {11'd 144,11'd 145};
    assign memory2[ 89] = {11'd 148,11'd 145};
    assign memory2[ 90] = {11'd 148,11'd 149};
    assign memory2[ 91] = {11'd 150,11'd 149};
    assign memory2[ 92] = {11'd 150,11'd 155};
    assign memory2[ 93] = {11'd 154,11'd 155};
    assign memory2[ 94] = {11'd 154,11'd 159};
    assign memory2[ 95] = {11'd 162,11'd 159};
    assign memory2[ 96] = {11'd 162,11'd 163};
    assign memory2[ 97] = {11'd 166,11'd 163};
    assign memory2[ 98] = {11'd 166,11'd 165};
    assign memory2[ 99] = {11'd 172,11'd 165};
    assign memory2[100] = {11'd 172,11'd 169};
    assign memory2[101] = {11'd 176,11'd 169};
    assign memory2[102] = {11'd 176,11'd 177};
    assign memory2[103] = {11'd 180,11'd 177};
    assign memory2[104] = {11'd 180,11'd 181};
    assign memory2[105] = {11'd 182,11'd 181};
    assign memory2[106] = {11'd 182,11'd 187};
    assign memory2[107] = {11'd 186,11'd 187};
    assign memory2[108] = {11'd 186,11'd 191};
    assign memory2[109] = {11'd 194,11'd 191};
    assign memory2[110] = {11'd 194,11'd 195};
    assign memory2[111] = {11'd 198,11'd 195};
    assign memory2[112] = {11'd 198,11'd 199};
    assign memory2[113] = {11'd 202,11'd 199};
    assign memory2[114] = {11'd 202,11'd 201};
    assign memory2[115] = {11'd 204,11'd 201};
    assign memory2[116] = {11'd 204,11'd 203};
    assign memory2[117] = {11'd 206,11'd 203};
    assign memory2[118] = {11'd 206,11'd 207};
    assign memory2[119] = {11'd 208,11'd 207};
    assign memory2[120] = {11'd 208,11'd 209};
    assign memory2[121] = {11'd 212,11'd 209};
    assign memory2[122] = {11'd 212,11'd 213};
    assign memory2[123] = {11'd 214,11'd 213};
    assign memory2[124] = {11'd 214,11'd 215};
    assign memory2[125] = {11'd 216,11'd 215};
    assign memory2[126] = {11'd 216,11'd 217};
    assign memory2[127] = {11'd 218,11'd 217};
    assign memory2[128] = {11'd 218,11'd 219};
    assign memory2[129] = {11'd 220,11'd 219};
    assign memory2[130] = {11'd 220,11'd 221};
    assign memory2[131] = {11'd 224,11'd 221};
    assign memory2[132] = {11'd 224,11'd 223};
    assign memory2[133] = {11'd 226,11'd 223};
    assign memory2[134] = {11'd 226,11'd 225};
    assign memory2[135] = {11'd 228,11'd 225};
    assign memory2[136] = {11'd 228,11'd 227};
    assign memory2[137] = {11'd 230,11'd 227};
    assign memory2[138] = {11'd 230,11'd 229};
    assign memory2[139] = {11'd 232,11'd 229};
    assign memory2[140] = {11'd 232,11'd 231};
    assign memory2[141] = {11'd 234,11'd 231};
    assign memory2[142] = {11'd 234,11'd 233};
    assign memory2[143] = {11'd 236,11'd 233};
    assign memory2[144] = {11'd 236,11'd 235};
    assign memory2[145] = {11'd 238,11'd 235};
    assign memory2[146] = {11'd 238,11'd 239};
    assign memory2[147] = {11'd 240,11'd 239};
    assign memory2[148] = {11'd 240,11'd 241};
    assign memory2[149] = {11'd 244,11'd 241};
    assign memory2[150] = {11'd 244,11'd 245};
    assign memory2[151] = {11'd 246,11'd 245};
    assign memory2[152] = {11'd 246,11'd 247};
    assign memory2[153] = {11'd 248,11'd 247};
    assign memory2[154] = {11'd 248,11'd 249};
    assign memory2[155] = {11'd 250,11'd 249};
    assign memory2[156] = {11'd 250,11'd 251};
    assign memory2[157] = {11'd 252,11'd 251};
    assign memory2[158] = {11'd 252,11'd 253};
    assign memory2[159] = {11'd 256,11'd 253};
    assign memory2[160] = {11'd 256,11'd 255};
    assign memory2[161] = {11'd 258,11'd 255};
    assign memory2[162] = {11'd 258,11'd 259};
    assign memory2[163] = {11'd 262,11'd 259};
    assign memory2[164] = {11'd 262,11'd 263};
    assign memory2[165] = {11'd 266,11'd 263};
    assign memory2[166] = {11'd 266,11'd 265};
    assign memory2[167] = {11'd 268,11'd 265};
    assign memory2[168] = {11'd 268,11'd 267};
    assign memory2[169] = {11'd 270,11'd 267};
    assign memory2[170] = {11'd 270,11'd 271};
    assign memory2[171] = {11'd 272,11'd 271};
    assign memory2[172] = {11'd 272,11'd 273};
    assign memory2[173] = {11'd 276,11'd 273};
    assign memory2[174] = {11'd 276,11'd 277};
    assign memory2[175] = {11'd 278,11'd 277};
    assign memory2[176] = {11'd 278,11'd 279};
    assign memory2[177] = {11'd 280,11'd 279};
    assign memory2[178] = {11'd 280,11'd 281};
    assign memory2[179] = {11'd 282,11'd 281};
    assign memory2[180] = {11'd 282,11'd 283};
    assign memory2[181] = {11'd 284,11'd 283};
    assign memory2[182] = {11'd 284,11'd 285};
    assign memory2[183] = {11'd 288,11'd 285};
    assign memory2[184] = {11'd 288,11'd 287};
    assign memory2[185] = {11'd 290,11'd 287};
    assign memory2[186] = {11'd 290,11'd 289};
    assign memory2[187] = {11'd 292,11'd 289};
    assign memory2[188] = {11'd 292,11'd 291};
    assign memory2[189] = {11'd 294,11'd 291};
    assign memory2[190] = {11'd 294,11'd 293};
    assign memory2[191] = {11'd 296,11'd 293};
    assign memory2[192] = {11'd 296,11'd 295};
    assign memory2[193] = {11'd 298,11'd 295};
    assign memory2[194] = {11'd 298,11'd 297};
    assign memory2[195] = {11'd 300,11'd 297};
    assign memory2[196] = {11'd 300,11'd 299};
    assign memory2[197] = {11'd 302,11'd 299};
    assign memory2[198] = {11'd 302,11'd 303};
    assign memory2[199] = {11'd 304,11'd 303};
    assign memory2[200] = {11'd 304,11'd 305};
    assign memory2[201] = {11'd 308,11'd 305};
    assign memory2[202] = {11'd 308,11'd 309};
    assign memory2[203] = {11'd 310,11'd 309};
    assign memory2[204] = {11'd 310,11'd 311};
    assign memory2[205] = {11'd 312,11'd 311};
    assign memory2[206] = {11'd 312,11'd 313};
    assign memory2[207] = {11'd 314,11'd 313};
    assign memory2[208] = {11'd 314,11'd 315};
    assign memory2[209] = {11'd 316,11'd 315};
    assign memory2[210] = {11'd 316,11'd 317};
    assign memory2[211] = {11'd 320,11'd 317};
    assign memory2[212] = {11'd 320,11'd 319};
    assign memory2[213] = {11'd 322,11'd 319};
    assign memory2[214] = {11'd 322,11'd 323};
    assign memory2[215] = {11'd 326,11'd 323};
    assign memory2[216] = {11'd 326,11'd 327};
    assign memory2[217] = {11'd 330,11'd 327};
    assign memory2[218] = {11'd 330,11'd 329};
    assign memory2[219] = {11'd 332,11'd 329};
    assign memory2[220] = {11'd 332,11'd 331};
    assign memory2[221] = {11'd 334,11'd 331};
    assign memory2[222] = {11'd 334,11'd 335};
    assign memory2[223] = {11'd 336,11'd 335};
    assign memory2[224] = {11'd 336,11'd 337};
    assign memory2[225] = {11'd 338,11'd 337};
    assign memory2[226] = {11'd 338,11'd 339};
    assign memory2[227] = {11'd 340,11'd 339};
    assign memory2[228] = {11'd 340,11'd 341};
    assign memory2[229] = {11'd 344,11'd 341};
    assign memory2[230] = {11'd 344,11'd 343};
    assign memory2[231] = {11'd 346,11'd 343};
    assign memory2[232] = {11'd 346,11'd 345};
    assign memory2[233] = {11'd 348,11'd 345};
    assign memory2[234] = {11'd 348,11'd 347};
    assign memory2[235] = {11'd 350,11'd 347};
    assign memory2[236] = {11'd 350,11'd 351};
    assign memory2[237] = {11'd 352,11'd 351};
    assign memory2[238] = {11'd 352,11'd 353};
    assign memory2[239] = {11'd 354,11'd 353};
    assign memory2[240] = {11'd 354,11'd 355};
    assign memory2[241] = {11'd 356,11'd 355};
    assign memory2[242] = {11'd 356,11'd 357};
    assign memory2[243] = {11'd 360,11'd 357};
    assign memory2[244] = {11'd 360,11'd 359};
    assign memory2[245] = {11'd 362,11'd 359};
    assign memory2[246] = {11'd 362,11'd 361};
    assign memory2[247] = {11'd 364,11'd 361};
    assign memory2[248] = {11'd 364,11'd 363};
    assign memory2[249] = {11'd 366,11'd 363};
    assign memory2[250] = {11'd 366,11'd 367};
    assign memory2[251] = {11'd 368,11'd 367};
    assign memory2[252] = {11'd 368,11'd 369};
    assign memory2[253] = {11'd 370,11'd 369};
    assign memory2[254] = {11'd 370,11'd 371};
    assign memory2[255] = {11'd 372,11'd 371};
    assign memory2[256] = {11'd 372,11'd 373};
    assign memory2[257] = {11'd 376,11'd 373};
    assign memory2[258] = {11'd 376,11'd 375};
    assign memory2[259] = {11'd 378,11'd 375};
    assign memory2[260] = {11'd 378,11'd 377};
    assign memory2[261] = {11'd 380,11'd 377};
    assign memory2[262] = {11'd 380,11'd 379};
    assign memory2[263] = {11'd 382,11'd 379};
    assign memory2[264] = {11'd 382,11'd 383};
    assign memory2[265] = {11'd 384,11'd 383};
    assign memory2[266] = {11'd 384,11'd 385};
    assign memory2[267] = {11'd 386,11'd 385};
    assign memory2[268] = {11'd 386,11'd 387};
    assign memory2[269] = {11'd 388,11'd 387};
    assign memory2[270] = {11'd 388,11'd 389};
    assign memory2[271] = {11'd 392,11'd 389};
    assign memory2[272] = {11'd 392,11'd 391};
    assign memory2[273] = {11'd 394,11'd 391};
    assign memory2[274] = {11'd 394,11'd 393};
    assign memory2[275] = {11'd 396,11'd 393};
    assign memory2[276] = {11'd 396,11'd 395};
    assign memory2[277] = {11'd 398,11'd 395};
    assign memory2[278] = {11'd 398,11'd 399};
    assign memory2[279] = {11'd 400,11'd 399};
    assign memory2[280] = {11'd 400,11'd 401};
    assign memory2[281] = {11'd 402,11'd 401};
    assign memory2[282] = {11'd 402,11'd 403};
    assign memory2[283] = {11'd 404,11'd 403};
    assign memory2[284] = {11'd 404,11'd 405};
    assign memory2[285] = {11'd 408,11'd 405};
    assign memory2[286] = {11'd 408,11'd 407};
    assign memory2[287] = {11'd 410,11'd 407};
    assign memory2[288] = {11'd 410,11'd 409};
    assign memory2[289] = {11'd 412,11'd 409};
    assign memory2[290] = {11'd 412,11'd 411};
    assign memory2[291] = {11'd 414,11'd 411};
    assign memory2[292] = {11'd 414,11'd 415};
    assign memory2[293] = {11'd 416,11'd 415};
    assign memory2[294] = {11'd 416,11'd 417};
    assign memory2[295] = {11'd 418,11'd 417};
    assign memory2[296] = {11'd 418,11'd 419};
    assign memory2[297] = {11'd 420,11'd 419};
    assign memory2[298] = {11'd 420,11'd 421};
    assign memory2[299] = {11'd 424,11'd 421};
    assign memory2[300] = {11'd 424,11'd 423};
    assign memory2[301] = {11'd 426,11'd 423};
    assign memory2[302] = {11'd 426,11'd 425};
    assign memory2[303] = {11'd 428,11'd 425};
    assign memory2[304] = {11'd 428,11'd 427};
    assign memory2[305] = {11'd 430,11'd 427};
    assign memory2[306] = {11'd 430,11'd 431};
    assign memory2[307] = {11'd 432,11'd 431};
    assign memory2[308] = {11'd 432,11'd 433};
    assign memory2[309] = {11'd 434,11'd 433};
    assign memory2[310] = {11'd 434,11'd 435};
    assign memory2[311] = {11'd 436,11'd 435};
    assign memory2[312] = {11'd 436,11'd 437};
    assign memory2[313] = {11'd 440,11'd 437};
    assign memory2[314] = {11'd 440,11'd 439};
    assign memory2[315] = {11'd 442,11'd 439};
    assign memory2[316] = {11'd 442,11'd 441};
    assign memory2[317] = {11'd 444,11'd 441};
    assign memory2[318] = {11'd 444,11'd 443};
    assign memory2[319] = {11'd 446,11'd 443};
    assign memory2[320] = {11'd 446,11'd 447};
    assign memory2[321] = {11'd 448,11'd 447};
    assign memory2[322] = {11'd 448,11'd 449};
    assign memory2[323] = {11'd 450,11'd 449};
    assign memory2[324] = {11'd 450,11'd 451};
    assign memory2[325] = {11'd 452,11'd 451};
    assign memory2[326] = {11'd 452,11'd 453};
    assign memory2[327] = {11'd 460,11'd 453};
    assign memory2[328] = {11'd 460,11'd 461};
    assign memory2[329] = {11'd 468,11'd 461};
    assign memory2[330] = {11'd 468,11'd 469};
    assign memory2[331] = {11'd 476,11'd 469};
    assign memory2[332] = {11'd 476,11'd 477};
    assign memory2[333] = {11'd 484,11'd 477};
    assign memory2[334] = {11'd 484,11'd 485};
    assign memory2[335] = {11'd 492,11'd 485};
    assign memory2[336] = {11'd 492,11'd 493};
    assign memory2[337] = {11'd 500,11'd 493};
    assign memory2[338] = {11'd 500,11'd 501};
    assign memory2[339] = {11'd 508,11'd 501};
    assign memory2[340] = {11'd 508,11'd 509};
    assign memory2[341] = {11'd 516,11'd 509};
    assign memory2[342] = {11'd 516,11'd 511};
    assign memory2[343] = {11'd 518,11'd 511};
    assign memory2[344] = {11'd 518,11'd 513};
    assign memory2[345] = {11'd 520,11'd 513};
    assign memory2[346] = {11'd 520,11'd 517};
    assign memory2[347] = {11'd 522,11'd 517};
    assign memory2[348] = {11'd 522,11'd 519};
    assign memory2[349] = {11'd 524,11'd 519};
    assign memory2[350] = {11'd 524,11'd 521};
    assign memory2[351] = {11'd 526,11'd 521};
    assign memory2[352] = {11'd 526,11'd 523};
    assign memory2[353] = {11'd 530,11'd 523};
    assign memory2[354] = {11'd 530,11'd 525};
    assign memory2[355] = {11'd 532,11'd 525};
    assign memory2[356] = {11'd 532,11'd 527};
    assign memory2[357] = {11'd 534,11'd 527};
    assign memory2[358] = {11'd 534,11'd 529};
    assign memory2[359] = {11'd 536,11'd 529};
    assign memory2[360] = {11'd 536,11'd 533};
    assign memory2[361] = {11'd 538,11'd 533};
    assign memory2[362] = {11'd 538,11'd 535};
    assign memory2[363] = {11'd 540,11'd 535};
    assign memory2[364] = {11'd 540,11'd 537};
    assign memory2[365] = {11'd 542,11'd 537};
    assign memory2[366] = {11'd 542,11'd 539};
    assign memory2[367] = {11'd 546,11'd 539};
    assign memory2[368] = {11'd 546,11'd 541};
    assign memory2[369] = {11'd 548,11'd 541};
    assign memory2[370] = {11'd 548,11'd 543};
    assign memory2[371] = {11'd 550,11'd 543};
    assign memory2[372] = {11'd 550,11'd 545};
    assign memory2[373] = {11'd 552,11'd 545};
    assign memory2[374] = {11'd 552,11'd 549};
    assign memory2[375] = {11'd 554,11'd 549};
    assign memory2[376] = {11'd 554,11'd 551};
    assign memory2[377] = {11'd 556,11'd 551};
    assign memory2[378] = {11'd 556,11'd 553};
    assign memory2[379] = {11'd 558,11'd 553};
    assign memory2[380] = {11'd 558,11'd 555};
    assign memory2[381] = {11'd 562,11'd 555};
    assign memory2[382] = {11'd 562,11'd 557};
    assign memory2[383] = {11'd 564,11'd 557};
    assign memory2[384] = {11'd 564,11'd 559};
    assign memory2[385] = {11'd 566,11'd 559};
    assign memory2[386] = {11'd 566,11'd 561};
    assign memory2[387] = {11'd 568,11'd 561};
    assign memory2[388] = {11'd 568,11'd 565};
    assign memory2[389] = {11'd 570,11'd 565};
    assign memory2[390] = {11'd 570,11'd 567};
    assign memory2[391] = {11'd 572,11'd 567};
    assign memory2[392] = {11'd 572,11'd 569};
    assign memory2[393] = {11'd 574,11'd 569};
    assign memory2[394] = {11'd 574,11'd 571};
    assign memory2[395] = {11'd 578,11'd 571};
    assign memory2[396] = {11'd 578,11'd 573};
    assign memory2[397] = {11'd 580,11'd 573};
    assign memory2[398] = {11'd 580,11'd 575};
    assign memory2[399] = {11'd 582,11'd 575};
    assign memory2[400] = {11'd 582,11'd 577};
    assign memory2[401] = {11'd 584,11'd 577};
    assign memory2[402] = {11'd 584,11'd 585};
    assign memory2[403] = {11'd 587,11'd 585};
    assign memory2[404] = {11'd 587,11'd 588};
    assign memory2[405] = {11'd 589,11'd 588};
    assign memory2[406] = {11'd 589,11'd 591};
    assign memory2[407] = {11'd 592,11'd 591};
    assign memory2[408] = {11'd 592,11'd 593};
    assign memory2[409] = {11'd 595,11'd 593};
    assign memory2[410] = {11'd 595,11'd 596};
    assign memory2[411] = {11'd 597,11'd 596};
    assign memory2[412] = {11'd 597,11'd 599};
    assign memory2[413] = {11'd 600,11'd 599};
    assign memory2[414] = {11'd 600,11'd 601};
    assign memory2[415] = {11'd 603,11'd 601};
    assign memory2[416] = {11'd 603,11'd 604};
    assign memory2[417] = {11'd 605,11'd 604};
    assign memory2[418] = {11'd 605,11'd 607};
    assign memory2[419] = {11'd 608,11'd 607};
    assign memory2[420] = {11'd 608,11'd 609};
    assign memory2[421] = {11'd 611,11'd 609};
    assign memory2[422] = {11'd 611,11'd 612};
    assign memory2[423] = {11'd 613,11'd 612};
    assign memory2[424] = {11'd 613,11'd 615};
    assign memory2[425] = {11'd 616,11'd 615};
    assign memory2[426] = {11'd 616,11'd 617};
    assign memory2[427] = {11'd 624,11'd 617};
    assign memory2[428] = {11'd 644,11'd 617};

    assign memory3[  0] = {11'd  10,11'd   7};
    assign memory3[  1] = {11'd  18,11'd   7};
    assign memory3[  2] = {11'd  18,11'd  15};
    assign memory3[  3] = {11'd  26,11'd  15};
    assign memory3[  4] = {11'd  26,11'd  17};
    assign memory3[  5] = {11'd  28,11'd  17};
    assign memory3[  6] = {11'd  28,11'd  21};
    assign memory3[  7] = {11'd  32,11'd  21};
    assign memory3[  8] = {11'd  32,11'd  25};
    assign memory3[  9] = {11'd  40,11'd  25};
    assign memory3[ 10] = {11'd  40,11'd  33};
    assign memory3[ 11] = {11'd  42,11'd  33};
    assign memory3[ 12] = {11'd  42,11'd  35};
    assign memory3[ 13] = {11'd  46,11'd  35};
    assign memory3[ 14] = {11'd  46,11'd  37};
    assign memory3[ 15] = {11'd  48,11'd  37};
    assign memory3[ 16] = {11'd  48,11'd  39};
    assign memory3[ 17] = {11'd  50,11'd  39};
    assign memory3[ 18] = {11'd  50,11'd  43};
    assign memory3[ 19] = {11'd  54,11'd  43};
    assign memory3[ 20] = {11'd  54,11'd  59};
    assign memory3[ 21] = {11'd  60,11'd  59};
    assign memory3[ 22] = {11'd  60,11'd  65};
    assign memory3[ 23] = {11'd  64,11'd  65};
    assign memory3[ 24] = {11'd  64,11'd  69};
    assign memory3[ 25] = {11'd  76,11'd  69};
    assign memory3[ 26] = {11'd  76,11'd  75};
    assign memory3[ 27] = {11'd  82,11'd  75};
    assign memory3[ 28] = {11'd  82,11'd  79};
    assign memory3[ 29] = {11'd  98,11'd  79};
    assign memory3[ 30] = {11'd  98,11'd  85};
    assign memory3[ 31] = {11'd 104,11'd  85};
    assign memory3[ 32] = {11'd 104,11'd  89};
    assign memory3[ 33] = {11'd 108,11'd  89};
    assign memory3[ 34] = {11'd 108,11'd 101};
    assign memory3[ 35] = {11'd 114,11'd 101};
    assign memory3[ 36] = {11'd 114,11'd 107};
    assign memory3[ 37] = {11'd 118,11'd 107};
    assign memory3[ 38] = {11'd 118,11'd 123};
    assign memory3[ 39] = {11'd 126,11'd 123};
    assign memory3[ 40] = {11'd 126,11'd 125};
    assign memory3[ 41] = {11'd 128,11'd 125};
    assign memory3[ 42] = {11'd 128,11'd 129};
    assign memory3[ 43] = {11'd 136,11'd 129};
    assign memory3[ 44] = {11'd 136,11'd 131};
    assign memory3[ 45] = {11'd 138,11'd 131};
    assign memory3[ 46] = {11'd 138,11'd 135};
    assign memory3[ 47] = {11'd 146,11'd 135};
    assign memory3[ 48] = {11'd 146,11'd 137};
    assign memory3[ 49] = {11'd 148,11'd 137};
    assign memory3[ 50] = {11'd 148,11'd 139};
    assign memory3[ 51] = {11'd 150,11'd 139};
    assign memory3[ 52] = {11'd 150,11'd 149};
    assign memory3[ 53] = {11'd 152,11'd 149};
    assign memory3[ 54] = {11'd 152,11'd 151};
    assign memory3[ 55] = {11'd 154,11'd 151};
    assign memory3[ 56] = {11'd 154,11'd 155};
    assign memory3[ 57] = {11'd 158,11'd 155};
    assign memory3[ 58] = {11'd 158,11'd 157};
    assign memory3[ 59] = {11'd 160,11'd 157};
    assign memory3[ 60] = {11'd 160,11'd 161};
    assign memory3[ 61] = {11'd 164,11'd 161};
    assign memory3[ 62] = {11'd 164,11'd 163};
    assign memory3[ 63] = {11'd 166,11'd 163};
    assign memory3[ 64] = {11'd 166,11'd 165};
    assign memory3[ 65] = {11'd 170,11'd 165};
    assign memory3[ 66] = {11'd 170,11'd 167};
    assign memory3[ 67] = {11'd 180,11'd 167};
    assign memory3[ 68] = {11'd 180,11'd 169};
    assign memory3[ 69] = {11'd 184,11'd 169};
    assign memory3[ 70] = {11'd 184,11'd 177};
    assign memory3[ 71] = {11'd 186,11'd 177};
    assign memory3[ 72] = {11'd 186,11'd 179};
    assign memory3[ 73] = {11'd 188,11'd 179};
    assign memory3[ 74] = {11'd 188,11'd 181};
    assign memory3[ 75] = {11'd 200,11'd 181};
    assign memory3[ 76] = {11'd 200,11'd 183};
    assign memory3[ 77] = {11'd 202,11'd 183};
    assign memory3[ 78] = {11'd 202,11'd 195};
    assign memory3[ 79] = {11'd 206,11'd 195};
    assign memory3[ 80] = {11'd 206,11'd 197};
    assign memory3[ 81] = {11'd 212,11'd 197};
    assign memory3[ 82] = {11'd 212,11'd 199};
    assign memory3[ 83] = {11'd 214,11'd 199};
    assign memory3[ 84] = {11'd 214,11'd 203};
    assign memory3[ 85] = {11'd 218,11'd 203};
    assign memory3[ 86] = {11'd 218,11'd 205};
    assign memory3[ 87] = {11'd 220,11'd 205};
    assign memory3[ 88] = {11'd 220,11'd 209};
    assign memory3[ 89] = {11'd 222,11'd 209};
    assign memory3[ 90] = {11'd 222,11'd 211};
    assign memory3[ 91] = {11'd 232,11'd 211};
    assign memory3[ 92] = {11'd 232,11'd 213};
    assign memory3[ 93] = {11'd 236,11'd 213};
    assign memory3[ 94] = {11'd 236,11'd 217};
    assign memory3[ 95] = {11'd 244,11'd 217};
    assign memory3[ 96] = {11'd 244,11'd 221};
    assign memory3[ 97] = {11'd 246,11'd 221};
    assign memory3[ 98] = {11'd 246,11'd 223};
    assign memory3[ 99] = {11'd 248,11'd 223};
    assign memory3[100] = {11'd 248,11'd 225};
    assign memory3[101] = {11'd 252,11'd 225};
    assign memory3[102] = {11'd 252,11'd 229};
    assign memory3[103] = {11'd 260,11'd 229};
    assign memory3[104] = {11'd 260,11'd 237};
    assign memory3[105] = {11'd 264,11'd 237};
    assign memory3[106] = {11'd 264,11'd 241};
    assign memory3[107] = {11'd 266,11'd 241};
    assign memory3[108] = {11'd 266,11'd 243};
    assign memory3[109] = {11'd 270,11'd 243};
    assign memory3[110] = {11'd 270,11'd 247};
    assign memory3[111] = {11'd 274,11'd 247};
    assign memory3[112] = {11'd 274,11'd 249};
    assign memory3[113] = {11'd 276,11'd 249};
    assign memory3[114] = {11'd 276,11'd 253};
    assign memory3[115] = {11'd 280,11'd 253};
    assign memory3[116] = {11'd 280,11'd 257};
    assign memory3[117] = {11'd 282,11'd 257};
    assign memory3[118] = {11'd 282,11'd 259};
    assign memory3[119] = {11'd 286,11'd 259};
    assign memory3[120] = {11'd 286,11'd 263};
    assign memory3[121] = {11'd 290,11'd 263};
    assign memory3[122] = {11'd 290,11'd 265};
    assign memory3[123] = {11'd 292,11'd 265};
    assign memory3[124] = {11'd 292,11'd 269};
    assign memory3[125] = {11'd 296,11'd 269};
    assign memory3[126] = {11'd 296,11'd 273};
    assign memory3[127] = {11'd 298,11'd 273};
    assign memory3[128] = {11'd 298,11'd 275};
    assign memory3[129] = {11'd 302,11'd 275};
    assign memory3[130] = {11'd 302,11'd 279};
    assign memory3[131] = {11'd 306,11'd 279};
    assign memory3[132] = {11'd 306,11'd 281};
    assign memory3[133] = {11'd 308,11'd 281};
    assign memory3[134] = {11'd 308,11'd 285};
    assign memory3[135] = {11'd 314,11'd 285};
    assign memory3[136] = {11'd 314,11'd 291};
    assign memory3[137] = {11'd 318,11'd 291};
    assign memory3[138] = {11'd 318,11'd 299};
    assign memory3[139] = {11'd 320,11'd 299};
    assign memory3[140] = {11'd 320,11'd 301};
    assign memory3[141] = {11'd 324,11'd 301};
    assign memory3[142] = {11'd 324,11'd 305};
    assign memory3[143] = {11'd 326,11'd 305};
    assign memory3[144] = {11'd 326,11'd 307};
    assign memory3[145] = {11'd 328,11'd 307};
    assign memory3[146] = {11'd 328,11'd 309};
    assign memory3[147] = {11'd 332,11'd 309};
    assign memory3[148] = {11'd 332,11'd 313};
    assign memory3[149] = {11'd 336,11'd 313};
    assign memory3[150] = {11'd 336,11'd 315};
    assign memory3[151] = {11'd 338,11'd 315};
    assign memory3[152] = {11'd 338,11'd 319};
    assign memory3[153] = {11'd 342,11'd 319};
    assign memory3[154] = {11'd 342,11'd 321};
    assign memory3[155] = {11'd 344,11'd 321};
    assign memory3[156] = {11'd 344,11'd 323};
    assign memory3[157] = {11'd 346,11'd 323};
    assign memory3[158] = {11'd 346,11'd 327};
    assign memory3[159] = {11'd 350,11'd 327};
    assign memory3[160] = {11'd 350,11'd 331};
    assign memory3[161] = {11'd 352,11'd 331};
    assign memory3[162] = {11'd 352,11'd 333};
    assign memory3[163] = {11'd 356,11'd 333};
    assign memory3[164] = {11'd 356,11'd 337};
    assign memory3[165] = {11'd 358,11'd 337};
    assign memory3[166] = {11'd 358,11'd 339};
    assign memory3[167] = {11'd 360,11'd 339};
    assign memory3[168] = {11'd 360,11'd 341};
    assign memory3[169] = {11'd 364,11'd 341};
    assign memory3[170] = {11'd 364,11'd 345};
    assign memory3[171] = {11'd 368,11'd 345};
    assign memory3[172] = {11'd 368,11'd 347};
    assign memory3[173] = {11'd 370,11'd 347};
    assign memory3[174] = {11'd 370,11'd 351};
    assign memory3[175] = {11'd 376,11'd 351};
    assign memory3[176] = {11'd 376,11'd 357};
    assign memory3[177] = {11'd 380,11'd 357};
    assign memory3[178] = {11'd 380,11'd 365};
    assign memory3[179] = {11'd 382,11'd 365};
    assign memory3[180] = {11'd 382,11'd 367};
    assign memory3[181] = {11'd 386,11'd 367};
    assign memory3[182] = {11'd 386,11'd 383};
    assign memory3[183] = {11'd 402,11'd 383};
    assign memory3[184] = {11'd 402,11'd 399};
    assign memory3[185] = {11'd 426,11'd 399};
    assign memory3[186] = {11'd 446,11'd 399};

    assign memory4[  0] = {11'd  10,11'd   7};
    assign memory4[  1] = {11'd  14,11'd   7};
    assign memory4[  2] = {11'd  14,11'd  15};
    assign memory4[  3] = {11'd  22,11'd  15};
    assign memory4[  4] = {11'd  22,11'd  17};
    assign memory4[  5] = {11'd  23,11'd  17};
    assign memory4[  6] = {11'd  23,11'd  20};
    assign memory4[  7] = {11'd  25,11'd  20};
    assign memory4[  8] = {11'd  25,11'd  28};
    assign memory4[  9] = {11'd  29,11'd  28};
    assign memory4[ 10] = {11'd  29,11'd  32};
    assign memory4[ 11] = {11'd  37,11'd  32};
    assign memory4[ 12] = {11'd  37,11'd  40};
    assign memory4[ 13] = {11'd  45,11'd  40};
    assign memory4[ 14] = {11'd  45,11'd  48};
    assign memory4[ 15] = {11'd  53,11'd  48};
    assign memory4[ 16] = {11'd  53,11'd  50};
    assign memory4[ 17] = {11'd  54,11'd  50};
    assign memory4[ 18] = {11'd  54,11'd  53};
    assign memory4[ 19] = {11'd  56,11'd  53};
    assign memory4[ 20] = {11'd  56,11'd  61};
    assign memory4[ 21] = {11'd  60,11'd  61};
    assign memory4[ 22] = {11'd  60,11'd  65};
    assign memory4[ 23] = {11'd  62,11'd  65};
    assign memory4[ 24] = {11'd  62,11'd  67};
    assign memory4[ 25] = {11'd  64,11'd  67};
    assign memory4[ 26] = {11'd  64,11'd  69};
    assign memory4[ 27] = {11'd  71,11'd  69};
    assign memory4[ 28] = {11'd  71,11'd  78};
    assign memory4[ 29] = {11'd  75,11'd  78};
    assign memory4[ 30] = {11'd  75,11'd  82};
    assign memory4[ 31] = {11'd  77,11'd  82};
    assign memory4[ 32] = {11'd  77,11'd  84};
    assign memory4[ 33] = {11'd  81,11'd  84};
    assign memory4[ 34] = {11'd  81,11'd  88};
    assign memory4[ 35] = {11'd  85,11'd  88};
    assign memory4[ 36] = {11'd  85,11'd  90};
    assign memory4[ 37] = {11'd  87,11'd  90};
    assign memory4[ 38] = {11'd  87,11'd  94};
    assign memory4[ 39] = {11'd  91,11'd  94};
    assign memory4[ 40] = {11'd  91,11'd  98};
    assign memory4[ 41] = {11'd  93,11'd  98};
    assign memory4[ 42] = {11'd  93,11'd 100};
    assign memory4[ 43] = {11'd  95,11'd 100};
    assign memory4[ 44] = {11'd  95,11'd 102};
    assign memory4[ 45] = {11'd  99,11'd 102};
    assign memory4[ 46] = {11'd  99,11'd 104};
    assign memory4[ 47] = {11'd 101,11'd 104};
    assign memory4[ 48] = {11'd 101,11'd 108};
    assign memory4[ 49] = {11'd 105,11'd 108};
    assign memory4[ 50] = {11'd 105,11'd 109};
    assign memory4[ 51] = {11'd 108,11'd 109};
    assign memory4[ 52] = {11'd 108,11'd 110};
    assign memory4[ 53] = {11'd 111,11'd 110};
    assign memory4[ 54] = {11'd 111,11'd 111};
    assign memory4[ 55] = {11'd 114,11'd 111};
    assign memory4[ 56] = {11'd 114,11'd 115};
    assign memory4[ 57] = {11'd 115,11'd 115};
    assign memory4[ 58] = {11'd 115,11'd 118};
    assign memory4[ 59] = {11'd 116,11'd 118};
    assign memory4[ 60] = {11'd 116,11'd 121};
    assign memory4[ 61] = {11'd 117,11'd 121};
    assign memory4[ 62] = {11'd 117,11'd 124};
    assign memory4[ 63] = {11'd 121,11'd 124};
    assign memory4[ 64] = {11'd 121,11'd 125};
    assign memory4[ 65] = {11'd 124,11'd 125};
    assign memory4[ 66] = {11'd 124,11'd 126};
    assign memory4[ 67] = {11'd 127,11'd 126};
    assign memory4[ 68] = {11'd 127,11'd 127};
    assign memory4[ 69] = {11'd 130,11'd 127};
    assign memory4[ 70] = {11'd 130,11'd 128};
    assign memory4[ 71] = {11'd 133,11'd 128};
    assign memory4[ 72] = {11'd 133,11'd 129};
    assign memory4[ 73] = {11'd 136,11'd 129};
    assign memory4[ 74] = {11'd 136,11'd 130};
    assign memory4[ 75] = {11'd 139,11'd 130};
    assign memory4[ 76] = {11'd 139,11'd 134};
    assign memory4[ 77] = {11'd 143,11'd 134};
    assign memory4[ 78] = {11'd 143,11'd 135};
    assign memory4[ 79] = {11'd 146,11'd 135};
    assign memory4[ 80] = {11'd 146,11'd 136};
    assign memory4[ 81] = {11'd 149,11'd 136};
    assign memory4[ 82] = {11'd 149,11'd 137};
    assign memory4[ 83] = {11'd 152,11'd 137};
    assign memory4[ 84] = {11'd 152,11'd 141};
    assign memory4[ 85] = {11'd 153,11'd 141};
    assign memory4[ 86] = {11'd 153,11'd 144};
    assign memory4[ 87] = {11'd 154,11'd 144};
    assign memory4[ 88] = {11'd 154,11'd 147};
    assign memory4[ 89] = {11'd 162,11'd 147};
    assign memory4[ 90] = {11'd 162,11'd 149};
    assign memory4[ 91] = {11'd 164,11'd 149};
    assign memory4[ 92] = {11'd 164,11'd 151};
    assign memory4[ 93] = {11'd 166,11'd 151};
    assign memory4[ 94] = {11'd 166,11'd 152};
    assign memory4[ 95] = {11'd 169,11'd 152};
    assign memory4[ 96] = {11'd 169,11'd 153};
    assign memory4[ 97] = {11'd 172,11'd 153};
    assign memory4[ 98] = {11'd 172,11'd 154};
    assign memory4[ 99] = {11'd 175,11'd 154};
    assign memory4[100] = {11'd 175,11'd 155};
    assign memory4[101] = {11'd 178,11'd 155};
    assign memory4[102] = {11'd 178,11'd 163};
    assign memory4[103] = {11'd 180,11'd 163};
    assign memory4[104] = {11'd 180,11'd 165};
    assign memory4[105] = {11'd 182,11'd 165};
    assign memory4[106] = {11'd 182,11'd 167};
    assign memory4[107] = {11'd 183,11'd 167};
    assign memory4[108] = {11'd 183,11'd 170};
    assign memory4[109] = {11'd 184,11'd 170};
    assign memory4[110] = {11'd 184,11'd 173};
    assign memory4[111] = {11'd 185,11'd 173};
    assign memory4[112] = {11'd 185,11'd 176};
    assign memory4[113] = {11'd 186,11'd 176};
    assign memory4[114] = {11'd 186,11'd 179};
    assign memory4[115] = {11'd 202,11'd 179};
    assign memory4[116] = {11'd 202,11'd 183};
    assign memory4[117] = {11'd 206,11'd 183};
    assign memory4[118] = {11'd 206,11'd 187};
    assign memory4[119] = {11'd 210,11'd 187};
    assign memory4[120] = {11'd 210,11'd 191};
    assign memory4[121] = {11'd 214,11'd 191};
    assign memory4[122] = {11'd 214,11'd 195};
    assign memory4[123] = {11'd 218,11'd 195};
    assign memory4[124] = {11'd 218,11'd 203};
    assign memory4[125] = {11'd 222,11'd 203};
    assign memory4[126] = {11'd 222,11'd 207};
    assign memory4[127] = {11'd 226,11'd 207};
    assign memory4[128] = {11'd 226,11'd 211};
    assign memory4[129] = {11'd 230,11'd 211};
    assign memory4[130] = {11'd 230,11'd 215};
    assign memory4[131] = {11'd 238,11'd 215};
    assign memory4[132] = {11'd 238,11'd 219};
    assign memory4[133] = {11'd 242,11'd 219};
    assign memory4[134] = {11'd 242,11'd 221};
    assign memory4[135] = {11'd 244,11'd 221};
    assign memory4[136] = {11'd 244,11'd 225};
    assign memory4[137] = {11'd 248,11'd 225};
    assign memory4[138] = {11'd 248,11'd 227};
    assign memory4[139] = {11'd 250,11'd 227};
    assign memory4[140] = {11'd 250,11'd 235};
    assign memory4[141] = {11'd 254,11'd 235};
    assign memory4[142] = {11'd 254,11'd 239};
    assign memory4[143] = {11'd 258,11'd 239};
    assign memory4[144] = {11'd 258,11'd 243};
    assign memory4[145] = {11'd 262,11'd 243};
    assign memory4[146] = {11'd 262,11'd 247};
    assign memory4[147] = {11'd 264,11'd 247};
    assign memory4[148] = {11'd 264,11'd 249};
    assign memory4[149] = {11'd 268,11'd 249};
    assign memory4[150] = {11'd 268,11'd 253};
    assign memory4[151] = {11'd 272,11'd 253};
    assign memory4[152] = {11'd 272,11'd 257};
    assign memory4[153] = {11'd 276,11'd 257};
    assign memory4[154] = {11'd 276,11'd 269};
    assign memory4[155] = {11'd 280,11'd 269};
    assign memory4[156] = {11'd 280,11'd 270};
    assign memory4[157] = {11'd 283,11'd 270};
    assign memory4[158] = {11'd 283,11'd 271};
    assign memory4[159] = {11'd 286,11'd 271};
    assign memory4[160] = {11'd 286,11'd 272};
    assign memory4[161] = {11'd 289,11'd 272};
    assign memory4[162] = {11'd 289,11'd 276};
    assign memory4[163] = {11'd 290,11'd 276};
    assign memory4[164] = {11'd 290,11'd 279};
    assign memory4[165] = {11'd 291,11'd 279};
    assign memory4[166] = {11'd 291,11'd 282};
    assign memory4[167] = {11'd 292,11'd 282};
    assign memory4[168] = {11'd 292,11'd 285};
    assign memory4[169] = {11'd 296,11'd 285};
    assign memory4[170] = {11'd 296,11'd 286};
    assign memory4[171] = {11'd 299,11'd 286};
    assign memory4[172] = {11'd 299,11'd 287};
    assign memory4[173] = {11'd 302,11'd 287};
    assign memory4[174] = {11'd 302,11'd 288};
    assign memory4[175] = {11'd 305,11'd 288};
    assign memory4[176] = {11'd 305,11'd 289};
    assign memory4[177] = {11'd 308,11'd 289};
    assign memory4[178] = {11'd 308,11'd 290};
    assign memory4[179] = {11'd 311,11'd 290};
    assign memory4[180] = {11'd 311,11'd 291};
    assign memory4[181] = {11'd 314,11'd 291};
    assign memory4[182] = {11'd 314,11'd 299};
    assign memory4[183] = {11'd 315,11'd 299};
    assign memory4[184] = {11'd 315,11'd 302};
    assign memory4[185] = {11'd 316,11'd 302};
    assign memory4[186] = {11'd 316,11'd 305};
    assign memory4[187] = {11'd 317,11'd 305};
    assign memory4[188] = {11'd 317,11'd 308};
    assign memory4[189] = {11'd 321,11'd 308};
    assign memory4[190] = {11'd 321,11'd 309};
    assign memory4[191] = {11'd 324,11'd 309};
    assign memory4[192] = {11'd 324,11'd 310};
    assign memory4[193] = {11'd 327,11'd 310};
    assign memory4[194] = {11'd 327,11'd 318};
    assign memory4[195] = {11'd 329,11'd 318};
    assign memory4[196] = {11'd 329,11'd 320};
    assign memory4[197] = {11'd 331,11'd 320};
    assign memory4[198] = {11'd 331,11'd 322};
    assign memory4[199] = {11'd 332,11'd 322};
    assign memory4[200] = {11'd 332,11'd 325};
    assign memory4[201] = {11'd 333,11'd 325};
    assign memory4[202] = {11'd 333,11'd 328};
    assign memory4[203] = {11'd 334,11'd 328};
    assign memory4[204] = {11'd 334,11'd 331};
    assign memory4[205] = {11'd 335,11'd 331};
    assign memory4[206] = {11'd 335,11'd 334};
    assign memory4[207] = {11'd 343,11'd 334};
    assign memory4[208] = {11'd 343,11'd 336};
    assign memory4[209] = {11'd 345,11'd 336};
    assign memory4[210] = {11'd 345,11'd 338};
    assign memory4[211] = {11'd 347,11'd 338};
    assign memory4[212] = {11'd 347,11'd 339};
    assign memory4[213] = {11'd 350,11'd 339};
    assign memory4[214] = {11'd 350,11'd 340};
    assign memory4[215] = {11'd 353,11'd 340};
    assign memory4[216] = {11'd 353,11'd 341};
    assign memory4[217] = {11'd 356,11'd 341};
    assign memory4[218] = {11'd 356,11'd 342};
    assign memory4[219] = {11'd 359,11'd 342};
    assign memory4[220] = {11'd 359,11'd 350};
    assign memory4[221] = {11'd 361,11'd 350};
    assign memory4[222] = {11'd 361,11'd 352};
    assign memory4[223] = {11'd 363,11'd 352};
    assign memory4[224] = {11'd 363,11'd 354};
    assign memory4[225] = {11'd 364,11'd 354};
    assign memory4[226] = {11'd 364,11'd 357};
    assign memory4[227] = {11'd 365,11'd 357};
    assign memory4[228] = {11'd 365,11'd 360};
    assign memory4[229] = {11'd 366,11'd 360};
    assign memory4[230] = {11'd 366,11'd 363};
    assign memory4[231] = {11'd 367,11'd 363};
    assign memory4[232] = {11'd 367,11'd 366};
    assign memory4[233] = {11'd 375,11'd 366};
    assign memory4[234] = {11'd 375,11'd 370};
    assign memory4[235] = {11'd 379,11'd 370};
    assign memory4[236] = {11'd 379,11'd 374};
    assign memory4[237] = {11'd 383,11'd 374};
    assign memory4[238] = {11'd 383,11'd 378};
    assign memory4[239] = {11'd 423,11'd 378};
    assign memory4[240] = {11'd 443,11'd 378};
    // ────────────────────────────────────────────────────────────────────────────────

endmodule
