//	How to use:	
//	1. Edit the songs on the Enter Song sheet.	
// 	2. Select this whole worksheet, copy it, and paste it into a new file.	
//	3. Save the file as song_rom.v.	

module drums_rom (
    input clk,						
	output reg [25:0] dout,						
	input [11:0] addr		
    );
        
    wire [25:0] memory [4095:0];  					
	always @(posedge clk)						
		dout = memory[addr];					

    parameter s1 = 538;
    parameter s2 = s1 + 529;
    parameter s3 = s2 + 411;

    assign memory[0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[1  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};
    assign memory[2  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[3  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[4  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[5  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[6  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[7  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[8  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[9  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[10 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[11 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[12 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[13 ] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[14 ] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[15 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[16 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[17 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[18 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[19 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[20 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[21 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[22 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[23 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[24 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[25 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[26 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[27 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[28 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[29 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[30 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[31 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[32 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[33 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[34 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[35 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[36 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[37 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[38 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[39 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[40 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[41 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[42 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[43 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[44 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[45 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[46 ] = {7'd7  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HKS
    assign memory[47 ] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[48 ] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[49 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[50 ] = {7'd5  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[51 ] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[52 ] = {7'd7  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSH
    assign memory[53 ] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[54 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[55 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[56 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[57 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[58 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[59 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[60 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[61 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[62 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[63 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[64 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[65 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[66 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[67 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[68 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[69 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[70 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[71 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[72 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[73 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[74 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[75 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[76 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[77 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[78 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[79 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[80 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[81 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[82 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[83 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[84 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[85 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[86 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[87 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[88 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[89 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[90 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[91 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[92 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[93 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[94 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[95 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[96 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[97 ] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[98 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[99 ] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[100] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[101] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[102] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[103] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[104] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[105] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[106] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[107] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[108] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[109] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[110] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[111] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[112] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[113] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[114] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[115] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[116] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[117] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[118] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[119] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[120] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[121] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[122] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[123] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[124] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[125] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[126] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[127] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[128] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[129] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[130] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[131] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[132] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[133] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[134] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[135] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[136] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[137] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[138] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[139] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[140] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[141] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[142] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[143] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[144] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[145] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[146] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[147] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[148] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[149] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[150] = {7'd5  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[151] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[152] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[153] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[154] = {7'd2  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[155] = {7'd5  , 8'd240, 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[156] = {7'd5  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KH
    assign memory[157] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[158] = {7'd2  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[159] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[160] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[161] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[162] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: KH
    assign memory[163] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[164] = {7'd5  , 8'd216, 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[165] = {7'd5  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KH
    assign memory[166] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[167] = {7'd2  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[168] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[169] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[170] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[171] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[172] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[173] = {7'd5  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KH
    assign memory[174] = {7'd5  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KH
    assign memory[175] = {7'd2  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[176] = {7'd1  , 8'd168, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[177] = {7'd4  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[178] = {7'd5  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KH
    assign memory[179] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[180] = {7'd2  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[181] = {7'd1  , 8'd120, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[182] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[183] = {7'd4  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[184] = {7'd5  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KH
    assign memory[185] = {7'd2  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[186] = {7'd1  , 8'd168, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[187] = {7'd4  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[188] = {7'd5  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KH
    assign memory[189] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[190] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[191] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[192] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[193] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[194] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[195] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[196] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[197] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[198] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[199] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[200] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[201] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[202] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[203] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[204] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[205] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[206] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[207] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[208] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[209] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[210] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[211] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[212] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[213] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[214] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[215] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[216] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[217] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[218] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[219] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[220] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[221] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[222] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[223] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[224] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[225] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[226] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[227] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[228] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[229] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[230] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[231] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[232] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[233] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[234] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[235] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[236] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[237] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[238] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[239] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[240] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[241] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[242] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[243] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[244] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[245] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[246] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[247] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[248] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[249] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[250] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[251] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[252] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[253] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[254] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[255] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[256] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[257] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[258] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[259] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[260] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[261] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[262] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[263] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[264] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[265] = {7'd1  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[266] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[267] = {7'd7  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSH
    assign memory[268] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[269] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[270] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[271] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[272] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[273] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[274] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[275] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[276] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[277] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[278] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[279] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[280] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[281] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[282] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[283] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[284] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[285] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[286] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[287] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[288] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[289] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[290] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[291] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[292] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[293] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[294] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[295] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[296] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[297] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[298] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[299] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[300] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[301] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[302] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[303] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[304] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[305] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[306] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[307] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[308] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[309] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[310] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[311] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[312] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[313] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[314] = {7'd1  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[315] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[316] = {7'd7  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSH
    assign memory[317] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[318] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[319] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[320] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[321] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[322] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[323] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[324] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[325] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[326] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[327] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[328] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[329] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[330] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[331] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[332] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[333] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[334] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[335] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[336] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[337] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[338] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[339] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[340] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[341] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[342] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[343] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[344] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[345] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[346] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[347] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[348] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[349] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[350] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[351] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[352] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[353] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[354] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[355] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[356] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[357] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[358] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[359] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[360] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[361] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[362] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[363] = {7'd1  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[364] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[365] = {7'd7  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSH
    assign memory[366] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[367] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[368] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[369] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[370] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[371] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[372] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[373] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[374] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[375] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[376] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[377] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[378] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[379] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[380] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[381] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[382] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[383] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[384] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[385] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[386] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[387] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[388] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[389] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[390] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[391] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[392] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[393] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[394] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[395] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[396] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[397] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[398] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[399] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[400] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[401] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[402] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[403] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[404] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[405] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[406] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[407] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[408] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[409] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[410] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[411] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[412] = {7'd1  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[413] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[414] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[415] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[416] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[417] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[418] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[419] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[420] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[421] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[422] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[423] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[424] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[425] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[426] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[427] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[428] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[429] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[430] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[431] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[432] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[433] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[434] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[435] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[436] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[437] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[438] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[439] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[440] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[441] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[442] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[443] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[444] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[445] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[446] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[447] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[448] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[449] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[450] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[451] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[452] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[453] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[454] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[455] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[456] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[457] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[458] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[459] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[460] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[461] = {7'd1  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[462] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[463] = {7'd7  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSH
    assign memory[464] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[465] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[466] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[467] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[468] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[469] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[470] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[471] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[472] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[473] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[474] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[475] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[476] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[477] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[478] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[479] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[480] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[481] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[482] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[483] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[484] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[485] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[486] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[487] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[488] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[489] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[490] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[491] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[492] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[493] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[494] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[495] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[496] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[497] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[498] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[499] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[500] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[501] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[502] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[503] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[504] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[505] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[506] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[507] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[508] = {7'd3  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[509] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[510] = {7'd1  , 8'd72 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[511] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[512] = {7'd7  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSH
    assign memory[513] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[514] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[515] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[516] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[517] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[518] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[519] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[520] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[521] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[522] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[523] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[524] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[525] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[526] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[527] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[528] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[529] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[530] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[531] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[532] = {7'd5  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HK
    assign memory[533] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[534] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[535] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[536] = {7'd0  , 8'd177, 7'd0  , 2'd0, 2'd0};
    assign memory[537] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song
    
    assign memory[s1+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s1+1  ] = {7'd10 , 8'd24 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+2  ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+3  ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+4  ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+5  ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+6  ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+7  ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+8  ] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+9  ] = {7'd6  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+10 ] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+11 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+12 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+13 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+14 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+15 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+16 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+17 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+18 ] = {7'd6  , 8'd60 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+19 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+20 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+21 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+22 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+23 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+24 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+25 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+26 ] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+27 ] = {7'd6  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+28 ] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+29 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+30 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+31 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+32 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+33 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+34 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+35 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+36 ] = {7'd6  , 8'd60 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+37 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+38 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+39 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+40 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+41 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+42 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+43 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+44 ] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+45 ] = {7'd6  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+46 ] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+47 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+48 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+49 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+50 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+51 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+52 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+53 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+54 ] = {7'd6  , 8'd60 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+55 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+56 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+57 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+58 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+59 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+60 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+61 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+62 ] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+63 ] = {7'd6  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+64 ] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+65 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+66 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+67 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+68 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+69 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+70 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+71 ] = {7'd10 , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: CS
    assign memory[s1+72 ] = {7'd2  , 8'd108, 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+73 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+74 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+75 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+76 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+77 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+78 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+79 ] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+80 ] = {7'd6  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+81 ] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+82 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+83 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+84 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+85 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+86 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+87 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+88 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+89 ] = {7'd6  , 8'd60 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+90 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+91 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+92 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+93 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+94 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+95 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+96 ] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+97 ] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+98 ] = {7'd6  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+99 ] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+100] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+101] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+102] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+103] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+104] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+105] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+106] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+107] = {7'd6  , 8'd60 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+108] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+109] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+110] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+111] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+112] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+113] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+114] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+115] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+116] = {7'd6  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+117] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+118] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+119] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+120] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+121] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+122] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+123] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+124] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+125] = {7'd6  , 8'd60 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+126] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+127] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+128] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+129] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+130] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+131] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+132] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+133] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+134] = {7'd6  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: HS
    assign memory[s1+135] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+136] = {7'd2  , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+137] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+138] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s1+139] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+140] = {7'd10 , 8'd36 , 7'd0  , 2'd0, 2'd0};   //note: SC
    assign memory[s1+141] = {7'd10 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: SC
    assign memory[s1+142] = {7'd14 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: SCH
    assign memory[s1+143] = {7'd10 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CS
    assign memory[s1+144] = {7'd10 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: SC
    assign memory[s1+145] = {7'd10 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: SC
    assign memory[s1+146] = {7'd11 , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+147] = {7'd3  , 8'd255, 7'd111, 2'd0, 2'd0};   //note: KS
    assign memory[s1+148] = {7'd0  , 8'd81 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+149] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+150] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+151] = {7'd3  , 8'd255, 7'd111, 2'd0, 2'd0};   //note: SK
    assign memory[s1+152] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+153] = {7'd3  , 8'd255, 7'd111, 2'd0, 2'd0};   //note: KS
    assign memory[s1+154] = {7'd0  , 8'd81 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+155] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+156] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+157] = {7'd3  , 8'd255, 7'd111, 2'd0, 2'd0};   //note: KS
    assign memory[s1+158] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+159] = {7'd3  , 8'd255, 7'd111, 2'd0, 2'd0};   //note: SK
    assign memory[s1+160] = {7'd0  , 8'd81 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+161] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+162] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+163] = {7'd3  , 8'd255, 7'd111, 2'd0, 2'd0};   //note: SK
    assign memory[s1+164] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+165] = {7'd3  , 8'd255, 7'd108, 2'd0, 2'd0};   //note: SK
    assign memory[s1+166] = {7'd0  , 8'd81 , 7'd0  , 2'd0, 2'd0};
    assign memory[s1+167] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+168] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+169] = {7'd11 , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: KCS
    assign memory[s1+170] = {7'd15 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: HKSC
    assign memory[s1+171] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: SCK
    assign memory[s1+172] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: KCS
    assign memory[s1+173] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+174] = {7'd11 , 8'd20 , 7'd0  , 2'd0, 2'd0};   //note: KCS
    assign memory[s1+175] = {7'd11 , 8'd44 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+176] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+177] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+178] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+179] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+180] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+181] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+182] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+183] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+184] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+185] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+186] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+187] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+188] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+189] = {7'd3  , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+190] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+191] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+192] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+193] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+194] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+195] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+196] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+197] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+198] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+199] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+200] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+201] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+202] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+203] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+204] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+205] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+206] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+207] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+208] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+209] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+210] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+211] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+212] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+213] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+214] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+215] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+216] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+217] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+218] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+219] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+220] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+221] = {7'd3  , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+222] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+223] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+224] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+225] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+226] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+227] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+228] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+229] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+230] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+231] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+232] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+233] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+234] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+235] = {7'd11 , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+236] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+237] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+238] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+239] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+240] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+241] = {7'd11 , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+242] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+243] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+244] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+245] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+246] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+247] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+248] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+249] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+250] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+251] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+252] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+253] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+254] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+255] = {7'd3  , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+256] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+257] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+258] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+259] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+260] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+261] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+262] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+263] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+264] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+265] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+266] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+267] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+268] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+269] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+270] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+271] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+272] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+273] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+274] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+275] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+276] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+277] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+278] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+279] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+280] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+281] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+282] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+283] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+284] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+285] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+286] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+287] = {7'd3  , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+288] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+289] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+290] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+291] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+292] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+293] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+294] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+295] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+296] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+297] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+298] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+299] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+300] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+301] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+302] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+303] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+304] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+305] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+306] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+307] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+308] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+309] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+310] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+311] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+312] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+313] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+314] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+315] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+316] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+317] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+318] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+319] = {7'd3  , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+320] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+321] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+322] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+323] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+324] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+325] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+326] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+327] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+328] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+329] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+330] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+331] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+332] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+333] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+334] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+335] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+336] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+337] = {7'd11 , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+338] = {7'd4  , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+339] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+340] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+341] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+342] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+343] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+344] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+345] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+346] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+347] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+348] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+349] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+350] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+351] = {7'd3  , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+352] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+353] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+354] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+355] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+356] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+357] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+358] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+359] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+360] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+361] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+362] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+363] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+364] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+365] = {7'd11 , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+366] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+367] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+368] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+369] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+370] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+371] = {7'd11 , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+372] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+373] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+374] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+375] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+376] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+377] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+378] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+379] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+380] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+381] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+382] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+383] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+384] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+385] = {7'd11 , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+386] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+387] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+388] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+389] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+390] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+391] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+392] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+393] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+394] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+395] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+396] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+397] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+398] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+399] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+400] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+401] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+402] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+403] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+404] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+405] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+406] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+407] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+408] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+409] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+410] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+411] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+412] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+413] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+414] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+415] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+416] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+417] = {7'd11 , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+418] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+419] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+420] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+421] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+422] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+423] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+424] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+425] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+426] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+427] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+428] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+429] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+430] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+431] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+432] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+433] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+434] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+435] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CKS
    assign memory[s1+436] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+437] = {7'd11 , 8'd32 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+438] = {7'd11 , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+439] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+440] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+441] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+442] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+443] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+444] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+445] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+446] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+447] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+448] = {7'd11 , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+449] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+450] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+451] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+452] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+453] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+454] = {7'd11 , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+455] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+456] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+457] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+458] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+459] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+460] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+461] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+462] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+463] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+464] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+465] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+466] = {7'd11 , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+467] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+468] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+469] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+470] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+471] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+472] = {7'd11 , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+473] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+474] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+475] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+476] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+477] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+478] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+479] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+480] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+481] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+482] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+483] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+484] = {7'd11 , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+485] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+486] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+487] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+488] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+489] = {7'd4  , 8'd56 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+490] = {7'd11 , 8'd40 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+491] = {7'd3  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+492] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+493] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+494] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KSC
    assign memory[s1+495] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+496] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+497] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+498] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: CSK
    assign memory[s1+499] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s1+500] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+501] = {7'd3  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s1+502] = {7'd11 , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+503] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+504] = {7'd11 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: SKC
    assign memory[s1+505] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s1+506] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s1+507] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+508] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+509] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+510] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+511] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+512] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+513] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+514] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+515] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+516] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+517] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+518] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+519] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+520] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+521] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+522] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+523] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+524] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+525] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+526] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+527] = {7'd0  , 8'd250, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+528] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s2+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s2+1  ] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+2  ] = {7'd0  , 8'd177, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+3  ] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};   //note: rest
    assign memory[s2+4  ] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+5  ] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+6  ] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};
    assign memory[s2+7  ] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};   //note: rest
    assign memory[s2+8  ] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+9  ] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+10 ] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};
    assign memory[s2+11 ] = {7'd8  , 8'd150, 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+12 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+13 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+14 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+15 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+16 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+17 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+18 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+19 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+20 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+21 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+22 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+23 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+24 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+25 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+26 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+27 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+28 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+29 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+30 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+31 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+32 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+33 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+34 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+35 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+36 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+37 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+38 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+39 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+40 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+41 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+42 ] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+43 ] = {7'd9  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: KC
    assign memory[s2+44 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+45 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+46 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+47 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+48 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+49 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+50 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+51 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+52 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+53 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+54 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+55 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+56 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+57 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+58 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+59 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+60 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+61 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+62 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+63 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+64 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+65 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+66 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+67 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+68 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+69 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+70 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+71 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+72 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+73 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+74 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+75 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+76 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+77 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+78 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+79 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+80 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+81 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+82 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+83 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+84 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+85 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+86 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+87 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+88 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+89 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+90 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+91 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+92 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+93 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+94 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+95 ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+96 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+97 ] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+98 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+99 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+100] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+101] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+102] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+103] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+104] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+105] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+106] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+107] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+108] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+109] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+110] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+111] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+112] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+113] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+114] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+115] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+116] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+117] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+118] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+119] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+120] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+121] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+122] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+123] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+124] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+125] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+126] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+127] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+128] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+129] = {7'd9  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s2+130] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+131] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+132] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+133] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+134] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+135] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+136] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+137] = {7'd10 , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: SC
    assign memory[s2+138] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+139] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+140] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+141] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+142] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+143] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+144] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+145] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+146] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+147] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+148] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+149] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+150] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+151] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+152] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+153] = {7'd8  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+154] = {7'd2  , 8'd255, 7'd97 , 2'd0, 2'd0};   //note: S
    assign memory[s2+155] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+156] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+157] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+158] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+159] = {7'd0  , 8'd255, 7'd97 , 2'd0, 2'd0};
    assign memory[s2+160] = {7'd0  , 8'd6  , 7'd0  , 2'd0, 2'd0};
    assign memory[s2+161] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+162] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+163] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+164] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+165] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+166] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+167] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+168] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+169] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+170] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+171] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+172] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+173] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+174] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+175] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+176] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+177] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+178] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+179] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+180] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+181] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+182] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+183] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+184] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+185] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+186] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+187] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+188] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+189] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+190] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+191] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+192] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+193] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+194] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+195] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+196] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+197] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+198] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+199] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+200] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+201] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+202] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+203] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+204] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+205] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+206] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+207] = {7'd2  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+208] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+209] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KC
    assign memory[s2+210] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+211] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+212] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+213] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+214] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+215] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+216] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+217] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+218] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+219] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+220] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+221] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+222] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+223] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+224] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+225] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+226] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s2+227] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+228] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+229] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+230] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+231] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+232] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+233] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+234] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+235] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+236] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+237] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+238] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+239] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+240] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+241] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+242] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+243] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KC
    assign memory[s2+244] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+245] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+246] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+247] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+248] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+249] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+250] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+251] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+252] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+253] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+254] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+255] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+256] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+257] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+258] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+259] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+260] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KC
    assign memory[s2+261] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+262] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+263] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+264] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+265] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+266] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+267] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+268] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+269] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+270] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+271] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+272] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+273] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+274] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+275] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+276] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+277] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s2+278] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+279] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+280] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+281] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+282] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+283] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+284] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+285] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+286] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+287] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+288] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+289] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+290] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+291] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+292] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+293] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+294] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s2+295] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+296] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+297] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+298] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+299] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+300] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+301] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+302] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+303] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+304] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+305] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+306] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+307] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+308] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+309] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+310] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+311] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s2+312] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+313] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+314] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+315] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+316] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+317] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+318] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+319] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+320] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+321] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+322] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+323] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+324] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+325] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+326] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+327] = {7'd2  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+328] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: KC
    assign memory[s2+329] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+330] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+331] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+332] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s2+333] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+334] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s2+335] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s2+336] = {7'd9  , 8'd30 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s2+337] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+338] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+339] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+340] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+341] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+342] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+343] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+344] = {7'd12 , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: CH
    assign memory[s2+345] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+346] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+347] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+348] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+349] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+350] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+351] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+352] = {7'd10 , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: CS
    assign memory[s2+353] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+354] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+355] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+356] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+357] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+358] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+359] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+360] = {7'd12 , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: HC
    assign memory[s2+361] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+362] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+363] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+364] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+365] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+366] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+367] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+368] = {7'd9  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s2+369] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+370] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+371] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+372] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+373] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+374] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+375] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+376] = {7'd12 , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: HC
    assign memory[s2+377] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+378] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+379] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+380] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+381] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+382] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+383] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+384] = {7'd10 , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: SC
    assign memory[s2+385] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+386] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+387] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+388] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+389] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+390] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+391] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+392] = {7'd10 , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: CS
    assign memory[s2+393] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+394] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+395] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+396] = {7'd10 , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: CS
    assign memory[s2+397] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+398] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+399] = {7'd8  , 8'd6  , 7'd0  , 2'd0, 2'd0};   //note: C
    assign memory[s2+400] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: KC
    assign memory[s2+401] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+402] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+403] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+404] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+405] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+406] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+407] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+408] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+409] = {7'd0  , 8'd154, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+410] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s3+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s3+1  ] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};
    assign memory[s3+2  ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+3  ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+4  ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+5  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+6  ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+7  ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+8  ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+9  ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+10 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+11 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+12 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+13 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+14 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+15 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+16 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+17 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+18 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+19 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+20 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+21 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+22 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+23 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+24 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+25 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+26 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+27 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+28 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+29 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+30 ] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+31 ] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+32 ] = {7'd2  , 8'd60 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+33 ] = {7'd2  , 8'd64 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+34 ] = {7'd3  , 8'd68 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s3+35 ] = {7'd1  , 8'd255, 7'd86 , 2'd0, 2'd0};   //note: K
    assign memory[s3+36 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+37 ] = {7'd2  , 8'd252, 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+38 ] = {7'd2  , 8'd64 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+39 ] = {7'd3  , 8'd68 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s3+40 ] = {7'd1  , 8'd255, 7'd86 , 2'd0, 2'd0};   //note: K
    assign memory[s3+41 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+42 ] = {7'd2  , 8'd252, 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+43 ] = {7'd2  , 8'd64 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+44 ] = {7'd3  , 8'd68 , 7'd0  , 2'd0, 2'd0};   //note: KS
    assign memory[s3+45 ] = {7'd1  , 8'd255, 7'd86 , 2'd0, 2'd0};   //note: K
    assign memory[s3+46 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+47 ] = {7'd2  , 8'd252, 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+48 ] = {7'd2  , 8'd64 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+49 ] = {7'd3  , 8'd68 , 7'd0  , 2'd0, 2'd0};   //note: SK
    assign memory[s3+50 ] = {7'd1  , 8'd255, 7'd86 , 2'd0, 2'd0};   //note: K
    assign memory[s3+51 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+52 ] = {7'd2  , 8'd60 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+53 ] = {7'd2  , 8'd64 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+54 ] = {7'd9  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s3+55 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+56 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+57 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+58 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+59 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+60 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+61 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+62 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+63 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+64 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+65 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+66 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+67 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+68 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+69 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+70 ] = {7'd9  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s3+71 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+72 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+73 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+74 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+75 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+76 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+77 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+78 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+79 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+80 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+81 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+82 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+83 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+84 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+85 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+86 ] = {7'd9  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s3+87 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+88 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+89 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+90 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+91 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+92 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+93 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+94 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+95 ] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+96 ] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+97 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+98 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+99 ] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+100] = {7'd12 , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: HC
    assign memory[s3+101] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+102] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+103] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+104] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+105] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+106] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+107] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+108] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+109] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+110] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+111] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+112] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+113] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+114] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+115] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+116] = {7'd12 , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: HC
    assign memory[s3+117] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+118] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+119] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+120] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+121] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+122] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+123] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+124] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+125] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+126] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+127] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+128] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+129] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+130] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+131] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+132] = {7'd12 , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: CH
    assign memory[s3+133] = {7'd1  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+134] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+135] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+136] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+137] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+138] = {7'd1  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+139] = {7'd4  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+140] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+141] = {7'd1  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+142] = {7'd4  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+143] = {7'd1  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+144] = {7'd4  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+145] = {7'd1  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+146] = {7'd4  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+147] = {7'd1  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+148] = {7'd4  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+149] = {7'd1  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+150] = {7'd4  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+151] = {7'd1  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+152] = {7'd4  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+153] = {7'd1  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+154] = {7'd4  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+155] = {7'd1  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+156] = {7'd4  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+157] = {7'd10 , 8'd255, 7'd86 , 2'd0, 2'd0};   //note: SC
    assign memory[s3+158] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+159] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+160] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+161] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+162] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+163] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+164] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+165] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+166] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+167] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+168] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+169] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+170] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+171] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+172] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+173] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+174] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+175] = {7'd0  , 8'd255, 7'd86 , 2'd0, 2'd0};
    assign memory[s3+176] = {7'd0  , 8'd3  , 7'd0  , 2'd0, 2'd0};
    assign memory[s3+177] = {7'd4  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+178] = {7'd1  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+179] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+180] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+181] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+182] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+183] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+184] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+185] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+186] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+187] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+188] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+189] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+190] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+191] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+192] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+193] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+194] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+195] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+196] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+197] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+198] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+199] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+200] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+201] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+202] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+203] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+204] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+205] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+206] = {7'd9  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: CK
    assign memory[s3+207] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+208] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+209] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+210] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+211] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+212] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+213] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+214] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+215] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+216] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+217] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+218] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+219] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+220] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+221] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+222] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+223] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+224] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+225] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+226] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+227] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+228] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+229] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+230] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+231] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+232] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+233] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+234] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+235] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+236] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+237] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+238] = {7'd9  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: KC
    assign memory[s3+239] = {7'd4  , 8'd144, 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+240] = {7'd2  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+241] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+242] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+243] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+244] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+245] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+246] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+247] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+248] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+249] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+250] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+251] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+252] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+253] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+254] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+255] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+256] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+257] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+258] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+259] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+260] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+261] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+262] = {7'd1  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: K
    assign memory[s3+263] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+264] = {7'd2  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: S
    assign memory[s3+265] = {7'd4  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: H
    assign memory[s3+266] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

endmodule							
