`timescale 1ns / 1ps

module hint_font_reader(
    input clk,
    input [4:0]character,
    input [9:0]x,
    input [4:0]y,
    output font_type
    );
    wire [12:0] hf_in;
    wire dout;
    hint_font_rom hfr(clk, hf_in, dout);
    
    assign hf_in = 12*character+x+348*y-12;
    assign font_type = (character==5'd0) ? 1'b0 : dout;
    
endmodule

module hint_font_rom(
    input clk,
    input [12:0] hf_in,
    output reg dout
    );
    wire memfont [6263:0];
    
    always @(posedge clk) begin
        dout = memfont[hf_in];
    end
    
    assign memfont[0   ] = 1'd0;
    assign memfont[1   ] = 1'd0;
    assign memfont[2   ] = 1'd0;
    assign memfont[3   ] = 1'd0;
    assign memfont[4   ] = 1'd0;
    assign memfont[5   ] = 1'd0;
    assign memfont[6   ] = 1'd0;
    assign memfont[7   ] = 1'd0;
    assign memfont[8   ] = 1'd0;
    assign memfont[9   ] = 1'd0;
    assign memfont[10  ] = 1'd0;
    assign memfont[11  ] = 1'd0;
    assign memfont[12  ] = 1'd0;
    assign memfont[13  ] = 1'd0;
    assign memfont[14  ] = 1'd0;
    assign memfont[15  ] = 1'd0;
    assign memfont[16  ] = 1'd0;
    assign memfont[17  ] = 1'd0;
    assign memfont[18  ] = 1'd0;
    assign memfont[19  ] = 1'd0;
    assign memfont[20  ] = 1'd0;
    assign memfont[21  ] = 1'd0;
    assign memfont[22  ] = 1'd0;
    assign memfont[23  ] = 1'd0;
    assign memfont[24  ] = 1'd0;
    assign memfont[25  ] = 1'd0;
    assign memfont[26  ] = 1'd0;
    assign memfont[27  ] = 1'd0;
    assign memfont[28  ] = 1'd0;
    assign memfont[29  ] = 1'd0;
    assign memfont[30  ] = 1'd0;
    assign memfont[31  ] = 1'd0;
    assign memfont[32  ] = 1'd0;
    assign memfont[33  ] = 1'd0;
    assign memfont[34  ] = 1'd0;
    assign memfont[35  ] = 1'd0;
    assign memfont[36  ] = 1'd0;
    assign memfont[37  ] = 1'd0;
    assign memfont[38  ] = 1'd0;
    assign memfont[39  ] = 1'd0;
    assign memfont[40  ] = 1'd0;
    assign memfont[41  ] = 1'd0;
    assign memfont[42  ] = 1'd0;
    assign memfont[43  ] = 1'd0;
    assign memfont[44  ] = 1'd0;
    assign memfont[45  ] = 1'd0;
    assign memfont[46  ] = 1'd0;
    assign memfont[47  ] = 1'd0;
    assign memfont[48  ] = 1'd0;
    assign memfont[49  ] = 1'd0;
    assign memfont[50  ] = 1'd0;
    assign memfont[51  ] = 1'd0;
    assign memfont[52  ] = 1'd0;
    assign memfont[53  ] = 1'd0;
    assign memfont[54  ] = 1'd0;
    assign memfont[55  ] = 1'd0;
    assign memfont[56  ] = 1'd0;
    assign memfont[57  ] = 1'd0;
    assign memfont[58  ] = 1'd0;
    assign memfont[59  ] = 1'd0;
    assign memfont[60  ] = 1'd0;
    assign memfont[61  ] = 1'd0;
    assign memfont[62  ] = 1'd0;
    assign memfont[63  ] = 1'd0;
    assign memfont[64  ] = 1'd0;
    assign memfont[65  ] = 1'd0;
    assign memfont[66  ] = 1'd0;
    assign memfont[67  ] = 1'd0;
    assign memfont[68  ] = 1'd0;
    assign memfont[69  ] = 1'd0;
    assign memfont[70  ] = 1'd0;
    assign memfont[71  ] = 1'd0;
    assign memfont[72  ] = 1'd0;
    assign memfont[73  ] = 1'd0;
    assign memfont[74  ] = 1'd0;
    assign memfont[75  ] = 1'd0;
    assign memfont[76  ] = 1'd0;
    assign memfont[77  ] = 1'd0;
    assign memfont[78  ] = 1'd0;
    assign memfont[79  ] = 1'd0;
    assign memfont[80  ] = 1'd0;
    assign memfont[81  ] = 1'd0;
    assign memfont[82  ] = 1'd0;
    assign memfont[83  ] = 1'd0;
    assign memfont[84  ] = 1'd0;
    assign memfont[85  ] = 1'd0;
    assign memfont[86  ] = 1'd0;
    assign memfont[87  ] = 1'd0;
    assign memfont[88  ] = 1'd0;
    assign memfont[89  ] = 1'd0;
    assign memfont[90  ] = 1'd0;
    assign memfont[91  ] = 1'd0;
    assign memfont[92  ] = 1'd0;
    assign memfont[93  ] = 1'd0;
    assign memfont[94  ] = 1'd0;
    assign memfont[95  ] = 1'd0;
    assign memfont[96  ] = 1'd0;
    assign memfont[97  ] = 1'd0;
    assign memfont[98  ] = 1'd0;
    assign memfont[99  ] = 1'd0;
    assign memfont[100 ] = 1'd0;
    assign memfont[101 ] = 1'd0;
    assign memfont[102 ] = 1'd0;
    assign memfont[103 ] = 1'd0;
    assign memfont[104 ] = 1'd0;
    assign memfont[105 ] = 1'd0;
    assign memfont[106 ] = 1'd0;
    assign memfont[107 ] = 1'd0;
    assign memfont[108 ] = 1'd0;
    assign memfont[109 ] = 1'd0;
    assign memfont[110 ] = 1'd0;
    assign memfont[111 ] = 1'd0;
    assign memfont[112 ] = 1'd0;
    assign memfont[113 ] = 1'd0;
    assign memfont[114 ] = 1'd0;
    assign memfont[115 ] = 1'd0;
    assign memfont[116 ] = 1'd0;
    assign memfont[117 ] = 1'd0;
    assign memfont[118 ] = 1'd0;
    assign memfont[119 ] = 1'd0;
    assign memfont[120 ] = 1'd0;
    assign memfont[121 ] = 1'd0;
    assign memfont[122 ] = 1'd0;
    assign memfont[123 ] = 1'd0;
    assign memfont[124 ] = 1'd0;
    assign memfont[125 ] = 1'd0;
    assign memfont[126 ] = 1'd0;
    assign memfont[127 ] = 1'd0;
    assign memfont[128 ] = 1'd0;
    assign memfont[129 ] = 1'd0;
    assign memfont[130 ] = 1'd0;
    assign memfont[131 ] = 1'd0;
    assign memfont[132 ] = 1'd0;
    assign memfont[133 ] = 1'd0;
    assign memfont[134 ] = 1'd0;
    assign memfont[135 ] = 1'd0;
    assign memfont[136 ] = 1'd0;
    assign memfont[137 ] = 1'd0;
    assign memfont[138 ] = 1'd0;
    assign memfont[139 ] = 1'd0;
    assign memfont[140 ] = 1'd0;
    assign memfont[141 ] = 1'd0;
    assign memfont[142 ] = 1'd0;
    assign memfont[143 ] = 1'd0;
    assign memfont[144 ] = 1'd0;
    assign memfont[145 ] = 1'd0;
    assign memfont[146 ] = 1'd0;
    assign memfont[147 ] = 1'd0;
    assign memfont[148 ] = 1'd0;
    assign memfont[149 ] = 1'd0;
    assign memfont[150 ] = 1'd0;
    assign memfont[151 ] = 1'd0;
    assign memfont[152 ] = 1'd0;
    assign memfont[153 ] = 1'd0;
    assign memfont[154 ] = 1'd0;
    assign memfont[155 ] = 1'd0;
    assign memfont[156 ] = 1'd0;
    assign memfont[157 ] = 1'd0;
    assign memfont[158 ] = 1'd0;
    assign memfont[159 ] = 1'd0;
    assign memfont[160 ] = 1'd0;
    assign memfont[161 ] = 1'd0;
    assign memfont[162 ] = 1'd0;
    assign memfont[163 ] = 1'd0;
    assign memfont[164 ] = 1'd0;
    assign memfont[165 ] = 1'd0;
    assign memfont[166 ] = 1'd0;
    assign memfont[167 ] = 1'd0;
    assign memfont[168 ] = 1'd0;
    assign memfont[169 ] = 1'd0;
    assign memfont[170 ] = 1'd0;
    assign memfont[171 ] = 1'd0;
    assign memfont[172 ] = 1'd0;
    assign memfont[173 ] = 1'd0;
    assign memfont[174 ] = 1'd0;
    assign memfont[175 ] = 1'd0;
    assign memfont[176 ] = 1'd0;
    assign memfont[177 ] = 1'd0;
    assign memfont[178 ] = 1'd0;
    assign memfont[179 ] = 1'd0;
    assign memfont[180 ] = 1'd0;
    assign memfont[181 ] = 1'd0;
    assign memfont[182 ] = 1'd0;
    assign memfont[183 ] = 1'd0;
    assign memfont[184 ] = 1'd0;
    assign memfont[185 ] = 1'd0;
    assign memfont[186 ] = 1'd0;
    assign memfont[187 ] = 1'd0;
    assign memfont[188 ] = 1'd0;
    assign memfont[189 ] = 1'd0;
    assign memfont[190 ] = 1'd0;
    assign memfont[191 ] = 1'd0;
    assign memfont[192 ] = 1'd0;
    assign memfont[193 ] = 1'd0;
    assign memfont[194 ] = 1'd0;
    assign memfont[195 ] = 1'd0;
    assign memfont[196 ] = 1'd0;
    assign memfont[197 ] = 1'd0;
    assign memfont[198 ] = 1'd0;
    assign memfont[199 ] = 1'd0;
    assign memfont[200 ] = 1'd0;
    assign memfont[201 ] = 1'd0;
    assign memfont[202 ] = 1'd0;
    assign memfont[203 ] = 1'd0;
    assign memfont[204 ] = 1'd0;
    assign memfont[205 ] = 1'd0;
    assign memfont[206 ] = 1'd0;
    assign memfont[207 ] = 1'd0;
    assign memfont[208 ] = 1'd0;
    assign memfont[209 ] = 1'd0;
    assign memfont[210 ] = 1'd0;
    assign memfont[211 ] = 1'd0;
    assign memfont[212 ] = 1'd0;
    assign memfont[213 ] = 1'd0;
    assign memfont[214 ] = 1'd0;
    assign memfont[215 ] = 1'd0;
    assign memfont[216 ] = 1'd0;
    assign memfont[217 ] = 1'd0;
    assign memfont[218 ] = 1'd0;
    assign memfont[219 ] = 1'd0;
    assign memfont[220 ] = 1'd0;
    assign memfont[221 ] = 1'd0;
    assign memfont[222 ] = 1'd0;
    assign memfont[223 ] = 1'd0;
    assign memfont[224 ] = 1'd0;
    assign memfont[225 ] = 1'd0;
    assign memfont[226 ] = 1'd0;
    assign memfont[227 ] = 1'd0;
    assign memfont[228 ] = 1'd0;
    assign memfont[229 ] = 1'd0;
    assign memfont[230 ] = 1'd0;
    assign memfont[231 ] = 1'd0;
    assign memfont[232 ] = 1'd0;
    assign memfont[233 ] = 1'd0;
    assign memfont[234 ] = 1'd0;
    assign memfont[235 ] = 1'd0;
    assign memfont[236 ] = 1'd0;
    assign memfont[237 ] = 1'd0;
    assign memfont[238 ] = 1'd0;
    assign memfont[239 ] = 1'd0;
    assign memfont[240 ] = 1'd0;
    assign memfont[241 ] = 1'd0;
    assign memfont[242 ] = 1'd0;
    assign memfont[243 ] = 1'd0;
    assign memfont[244 ] = 1'd0;
    assign memfont[245 ] = 1'd0;
    assign memfont[246 ] = 1'd0;
    assign memfont[247 ] = 1'd0;
    assign memfont[248 ] = 1'd0;
    assign memfont[249 ] = 1'd0;
    assign memfont[250 ] = 1'd0;
    assign memfont[251 ] = 1'd0;
    assign memfont[252 ] = 1'd0;
    assign memfont[253 ] = 1'd0;
    assign memfont[254 ] = 1'd0;
    assign memfont[255 ] = 1'd0;
    assign memfont[256 ] = 1'd0;
    assign memfont[257 ] = 1'd0;
    assign memfont[258 ] = 1'd0;
    assign memfont[259 ] = 1'd0;
    assign memfont[260 ] = 1'd0;
    assign memfont[261 ] = 1'd0;
    assign memfont[262 ] = 1'd0;
    assign memfont[263 ] = 1'd0;
    assign memfont[264 ] = 1'd0;
    assign memfont[265 ] = 1'd0;
    assign memfont[266 ] = 1'd0;
    assign memfont[267 ] = 1'd0;
    assign memfont[268 ] = 1'd0;
    assign memfont[269 ] = 1'd0;
    assign memfont[270 ] = 1'd0;
    assign memfont[271 ] = 1'd0;
    assign memfont[272 ] = 1'd0;
    assign memfont[273 ] = 1'd0;
    assign memfont[274 ] = 1'd0;
    assign memfont[275 ] = 1'd0;
    assign memfont[276 ] = 1'd0;
    assign memfont[277 ] = 1'd0;
    assign memfont[278 ] = 1'd0;
    assign memfont[279 ] = 1'd0;
    assign memfont[280 ] = 1'd0;
    assign memfont[281 ] = 1'd0;
    assign memfont[282 ] = 1'd0;
    assign memfont[283 ] = 1'd0;
    assign memfont[284 ] = 1'd0;
    assign memfont[285 ] = 1'd0;
    assign memfont[286 ] = 1'd0;
    assign memfont[287 ] = 1'd0;
    assign memfont[288 ] = 1'd0;
    assign memfont[289 ] = 1'd0;
    assign memfont[290 ] = 1'd0;
    assign memfont[291 ] = 1'd0;
    assign memfont[292 ] = 1'd0;
    assign memfont[293 ] = 1'd0;
    assign memfont[294 ] = 1'd0;
    assign memfont[295 ] = 1'd0;
    assign memfont[296 ] = 1'd0;
    assign memfont[297 ] = 1'd0;
    assign memfont[298 ] = 1'd0;
    assign memfont[299 ] = 1'd0;
    assign memfont[300 ] = 1'd0;
    assign memfont[301 ] = 1'd0;
    assign memfont[302 ] = 1'd0;
    assign memfont[303 ] = 1'd0;
    assign memfont[304 ] = 1'd0;
    assign memfont[305 ] = 1'd0;
    assign memfont[306 ] = 1'd0;
    assign memfont[307 ] = 1'd0;
    assign memfont[308 ] = 1'd0;
    assign memfont[309 ] = 1'd0;
    assign memfont[310 ] = 1'd0;
    assign memfont[311 ] = 1'd0;
    assign memfont[312 ] = 1'd0;
    assign memfont[313 ] = 1'd0;
    assign memfont[314 ] = 1'd0;
    assign memfont[315 ] = 1'd0;
    assign memfont[316 ] = 1'd0;
    assign memfont[317 ] = 1'd1;
    assign memfont[318 ] = 1'd1;
    assign memfont[319 ] = 1'd0;
    assign memfont[320 ] = 1'd0;
    assign memfont[321 ] = 1'd0;
    assign memfont[322 ] = 1'd0;
    assign memfont[323 ] = 1'd0;
    assign memfont[324 ] = 1'd0;
    assign memfont[325 ] = 1'd0;
    assign memfont[326 ] = 1'd0;
    assign memfont[327 ] = 1'd0;
    assign memfont[328 ] = 1'd0;
    assign memfont[329 ] = 1'd0;
    assign memfont[330 ] = 1'd0;
    assign memfont[331 ] = 1'd0;
    assign memfont[332 ] = 1'd0;
    assign memfont[333 ] = 1'd0;
    assign memfont[334 ] = 1'd0;
    assign memfont[335 ] = 1'd0;
    assign memfont[336 ] = 1'd0;
    assign memfont[337 ] = 1'd0;
    assign memfont[338 ] = 1'd0;
    assign memfont[339 ] = 1'd0;
    assign memfont[340 ] = 1'd0;
    assign memfont[341 ] = 1'd0;
    assign memfont[342 ] = 1'd0;
    assign memfont[343 ] = 1'd0;
    assign memfont[344 ] = 1'd0;
    assign memfont[345 ] = 1'd0;
    assign memfont[346 ] = 1'd0;
    assign memfont[347 ] = 1'd0;
    assign memfont[348 ] = 1'd0;
    assign memfont[349 ] = 1'd0;
    assign memfont[350 ] = 1'd0;
    assign memfont[351 ] = 1'd0;
    assign memfont[352 ] = 1'd0;
    assign memfont[353 ] = 1'd1;
    assign memfont[354 ] = 1'd1;
    assign memfont[355 ] = 1'd0;
    assign memfont[356 ] = 1'd0;
    assign memfont[357 ] = 1'd0;
    assign memfont[358 ] = 1'd0;
    assign memfont[359 ] = 1'd0;
    assign memfont[360 ] = 1'd0;
    assign memfont[361 ] = 1'd1;
    assign memfont[362 ] = 1'd1;
    assign memfont[363 ] = 1'd1;
    assign memfont[364 ] = 1'd1;
    assign memfont[365 ] = 1'd1;
    assign memfont[366 ] = 1'd0;
    assign memfont[367 ] = 1'd0;
    assign memfont[368 ] = 1'd0;
    assign memfont[369 ] = 1'd0;
    assign memfont[370 ] = 1'd0;
    assign memfont[371 ] = 1'd0;
    assign memfont[372 ] = 1'd0;
    assign memfont[373 ] = 1'd0;
    assign memfont[374 ] = 1'd0;
    assign memfont[375 ] = 1'd0;
    assign memfont[376 ] = 1'd0;
    assign memfont[377 ] = 1'd1;
    assign memfont[378 ] = 1'd1;
    assign memfont[379 ] = 1'd1;
    assign memfont[380 ] = 1'd0;
    assign memfont[381 ] = 1'd0;
    assign memfont[382 ] = 1'd0;
    assign memfont[383 ] = 1'd0;
    assign memfont[384 ] = 1'd0;
    assign memfont[385 ] = 1'd1;
    assign memfont[386 ] = 1'd1;
    assign memfont[387 ] = 1'd1;
    assign memfont[388 ] = 1'd0;
    assign memfont[389 ] = 1'd0;
    assign memfont[390 ] = 1'd0;
    assign memfont[391 ] = 1'd0;
    assign memfont[392 ] = 1'd0;
    assign memfont[393 ] = 1'd0;
    assign memfont[394 ] = 1'd0;
    assign memfont[395 ] = 1'd0;
    assign memfont[396 ] = 1'd0;
    assign memfont[397 ] = 1'd1;
    assign memfont[398 ] = 1'd1;
    assign memfont[399 ] = 1'd1;
    assign memfont[400 ] = 1'd1;
    assign memfont[401 ] = 1'd1;
    assign memfont[402 ] = 1'd1;
    assign memfont[403 ] = 1'd1;
    assign memfont[404 ] = 1'd1;
    assign memfont[405 ] = 1'd1;
    assign memfont[406 ] = 1'd0;
    assign memfont[407 ] = 1'd0;
    assign memfont[408 ] = 1'd0;
    assign memfont[409 ] = 1'd1;
    assign memfont[410 ] = 1'd1;
    assign memfont[411 ] = 1'd1;
    assign memfont[412 ] = 1'd1;
    assign memfont[413 ] = 1'd1;
    assign memfont[414 ] = 1'd1;
    assign memfont[415 ] = 1'd1;
    assign memfont[416 ] = 1'd1;
    assign memfont[417 ] = 1'd1;
    assign memfont[418 ] = 1'd1;
    assign memfont[419 ] = 1'd0;
    assign memfont[420 ] = 1'd0;
    assign memfont[421 ] = 1'd0;
    assign memfont[422 ] = 1'd0;
    assign memfont[423 ] = 1'd0;
    assign memfont[424 ] = 1'd0;
    assign memfont[425 ] = 1'd1;
    assign memfont[426 ] = 1'd1;
    assign memfont[427 ] = 1'd0;
    assign memfont[428 ] = 1'd0;
    assign memfont[429 ] = 1'd0;
    assign memfont[430 ] = 1'd0;
    assign memfont[431 ] = 1'd0;
    assign memfont[432 ] = 1'd0;
    assign memfont[433 ] = 1'd1;
    assign memfont[434 ] = 1'd1;
    assign memfont[435 ] = 1'd0;
    assign memfont[436 ] = 1'd0;
    assign memfont[437 ] = 1'd0;
    assign memfont[438 ] = 1'd0;
    assign memfont[439 ] = 1'd0;
    assign memfont[440 ] = 1'd0;
    assign memfont[441 ] = 1'd1;
    assign memfont[442 ] = 1'd1;
    assign memfont[443 ] = 1'd0;
    assign memfont[444 ] = 1'd0;
    assign memfont[445 ] = 1'd0;
    assign memfont[446 ] = 1'd0;
    assign memfont[447 ] = 1'd0;
    assign memfont[448 ] = 1'd0;
    assign memfont[449 ] = 1'd1;
    assign memfont[450 ] = 1'd1;
    assign memfont[451 ] = 1'd0;
    assign memfont[452 ] = 1'd0;
    assign memfont[453 ] = 1'd0;
    assign memfont[454 ] = 1'd0;
    assign memfont[455 ] = 1'd0;
    assign memfont[456 ] = 1'd0;
    assign memfont[457 ] = 1'd0;
    assign memfont[458 ] = 1'd0;
    assign memfont[459 ] = 1'd0;
    assign memfont[460 ] = 1'd0;
    assign memfont[461 ] = 1'd0;
    assign memfont[462 ] = 1'd0;
    assign memfont[463 ] = 1'd0;
    assign memfont[464 ] = 1'd1;
    assign memfont[465 ] = 1'd1;
    assign memfont[466 ] = 1'd1;
    assign memfont[467 ] = 1'd0;
    assign memfont[468 ] = 1'd0;
    assign memfont[469 ] = 1'd1;
    assign memfont[470 ] = 1'd1;
    assign memfont[471 ] = 1'd0;
    assign memfont[472 ] = 1'd0;
    assign memfont[473 ] = 1'd0;
    assign memfont[474 ] = 1'd0;
    assign memfont[475 ] = 1'd0;
    assign memfont[476 ] = 1'd0;
    assign memfont[477 ] = 1'd1;
    assign memfont[478 ] = 1'd1;
    assign memfont[479 ] = 1'd0;
    assign memfont[480 ] = 1'd0;
    assign memfont[481 ] = 1'd1;
    assign memfont[482 ] = 1'd1;
    assign memfont[483 ] = 1'd0;
    assign memfont[484 ] = 1'd0;
    assign memfont[485 ] = 1'd0;
    assign memfont[486 ] = 1'd0;
    assign memfont[487 ] = 1'd0;
    assign memfont[488 ] = 1'd0;
    assign memfont[489 ] = 1'd0;
    assign memfont[490 ] = 1'd0;
    assign memfont[491 ] = 1'd0;
    assign memfont[492 ] = 1'd0;
    assign memfont[493 ] = 1'd1;
    assign memfont[494 ] = 1'd1;
    assign memfont[495 ] = 1'd1;
    assign memfont[496 ] = 1'd0;
    assign memfont[497 ] = 1'd0;
    assign memfont[498 ] = 1'd0;
    assign memfont[499 ] = 1'd0;
    assign memfont[500 ] = 1'd1;
    assign memfont[501 ] = 1'd1;
    assign memfont[502 ] = 1'd1;
    assign memfont[503 ] = 1'd0;
    assign memfont[504 ] = 1'd0;
    assign memfont[505 ] = 1'd1;
    assign memfont[506 ] = 1'd1;
    assign memfont[507 ] = 1'd0;
    assign memfont[508 ] = 1'd0;
    assign memfont[509 ] = 1'd0;
    assign memfont[510 ] = 1'd0;
    assign memfont[511 ] = 1'd0;
    assign memfont[512 ] = 1'd0;
    assign memfont[513 ] = 1'd1;
    assign memfont[514 ] = 1'd1;
    assign memfont[515 ] = 1'd0;
    assign memfont[516 ] = 1'd0;
    assign memfont[517 ] = 1'd0;
    assign memfont[518 ] = 1'd0;
    assign memfont[519 ] = 1'd0;
    assign memfont[520 ] = 1'd1;
    assign memfont[521 ] = 1'd1;
    assign memfont[522 ] = 1'd1;
    assign memfont[523 ] = 1'd0;
    assign memfont[524 ] = 1'd0;
    assign memfont[525 ] = 1'd0;
    assign memfont[526 ] = 1'd0;
    assign memfont[527 ] = 1'd0;
    assign memfont[528 ] = 1'd0;
    assign memfont[529 ] = 1'd1;
    assign memfont[530 ] = 1'd1;
    assign memfont[531 ] = 1'd1;
    assign memfont[532 ] = 1'd1;
    assign memfont[533 ] = 1'd1;
    assign memfont[534 ] = 1'd0;
    assign memfont[535 ] = 1'd0;
    assign memfont[536 ] = 1'd0;
    assign memfont[537 ] = 1'd0;
    assign memfont[538 ] = 1'd0;
    assign memfont[539 ] = 1'd0;
    assign memfont[540 ] = 1'd0;
    assign memfont[541 ] = 1'd0;
    assign memfont[542 ] = 1'd0;
    assign memfont[543 ] = 1'd0;
    assign memfont[544 ] = 1'd1;
    assign memfont[545 ] = 1'd1;
    assign memfont[546 ] = 1'd1;
    assign memfont[547 ] = 1'd0;
    assign memfont[548 ] = 1'd0;
    assign memfont[549 ] = 1'd0;
    assign memfont[550 ] = 1'd0;
    assign memfont[551 ] = 1'd0;
    assign memfont[552 ] = 1'd0;
    assign memfont[553 ] = 1'd1;
    assign memfont[554 ] = 1'd1;
    assign memfont[555 ] = 1'd1;
    assign memfont[556 ] = 1'd1;
    assign memfont[557 ] = 1'd1;
    assign memfont[558 ] = 1'd0;
    assign memfont[559 ] = 1'd0;
    assign memfont[560 ] = 1'd0;
    assign memfont[561 ] = 1'd0;
    assign memfont[562 ] = 1'd0;
    assign memfont[563 ] = 1'd0;
    assign memfont[564 ] = 1'd0;
    assign memfont[565 ] = 1'd0;
    assign memfont[566 ] = 1'd0;
    assign memfont[567 ] = 1'd0;
    assign memfont[568 ] = 1'd1;
    assign memfont[569 ] = 1'd1;
    assign memfont[570 ] = 1'd1;
    assign memfont[571 ] = 1'd0;
    assign memfont[572 ] = 1'd0;
    assign memfont[573 ] = 1'd0;
    assign memfont[574 ] = 1'd0;
    assign memfont[575 ] = 1'd0;
    assign memfont[576 ] = 1'd0;
    assign memfont[577 ] = 1'd1;
    assign memfont[578 ] = 1'd1;
    assign memfont[579 ] = 1'd1;
    assign memfont[580 ] = 1'd1;
    assign memfont[581 ] = 1'd1;
    assign memfont[582 ] = 1'd1;
    assign memfont[583 ] = 1'd1;
    assign memfont[584 ] = 1'd1;
    assign memfont[585 ] = 1'd1;
    assign memfont[586 ] = 1'd1;
    assign memfont[587 ] = 1'd0;
    assign memfont[588 ] = 1'd0;
    assign memfont[589 ] = 1'd1;
    assign memfont[590 ] = 1'd1;
    assign memfont[591 ] = 1'd0;
    assign memfont[592 ] = 1'd0;
    assign memfont[593 ] = 1'd0;
    assign memfont[594 ] = 1'd0;
    assign memfont[595 ] = 1'd0;
    assign memfont[596 ] = 1'd0;
    assign memfont[597 ] = 1'd1;
    assign memfont[598 ] = 1'd1;
    assign memfont[599 ] = 1'd0;
    assign memfont[600 ] = 1'd1;
    assign memfont[601 ] = 1'd1;
    assign memfont[602 ] = 1'd0;
    assign memfont[603 ] = 1'd0;
    assign memfont[604 ] = 1'd0;
    assign memfont[605 ] = 1'd0;
    assign memfont[606 ] = 1'd0;
    assign memfont[607 ] = 1'd0;
    assign memfont[608 ] = 1'd0;
    assign memfont[609 ] = 1'd1;
    assign memfont[610 ] = 1'd1;
    assign memfont[611 ] = 1'd0;
    assign memfont[612 ] = 1'd1;
    assign memfont[613 ] = 1'd1;
    assign memfont[614 ] = 1'd0;
    assign memfont[615 ] = 1'd0;
    assign memfont[616 ] = 1'd0;
    assign memfont[617 ] = 1'd1;
    assign memfont[618 ] = 1'd1;
    assign memfont[619 ] = 1'd0;
    assign memfont[620 ] = 1'd0;
    assign memfont[621 ] = 1'd1;
    assign memfont[622 ] = 1'd1;
    assign memfont[623 ] = 1'd1;
    assign memfont[624 ] = 1'd0;
    assign memfont[625 ] = 1'd1;
    assign memfont[626 ] = 1'd1;
    assign memfont[627 ] = 1'd0;
    assign memfont[628 ] = 1'd0;
    assign memfont[629 ] = 1'd0;
    assign memfont[630 ] = 1'd0;
    assign memfont[631 ] = 1'd0;
    assign memfont[632 ] = 1'd0;
    assign memfont[633 ] = 1'd1;
    assign memfont[634 ] = 1'd1;
    assign memfont[635 ] = 1'd0;
    assign memfont[636 ] = 1'd1;
    assign memfont[637 ] = 1'd1;
    assign memfont[638 ] = 1'd1;
    assign memfont[639 ] = 1'd0;
    assign memfont[640 ] = 1'd0;
    assign memfont[641 ] = 1'd0;
    assign memfont[642 ] = 1'd0;
    assign memfont[643 ] = 1'd0;
    assign memfont[644 ] = 1'd0;
    assign memfont[645 ] = 1'd1;
    assign memfont[646 ] = 1'd1;
    assign memfont[647 ] = 1'd0;
    assign memfont[648 ] = 1'd0;
    assign memfont[649 ] = 1'd1;
    assign memfont[650 ] = 1'd1;
    assign memfont[651 ] = 1'd1;
    assign memfont[652 ] = 1'd1;
    assign memfont[653 ] = 1'd1;
    assign memfont[654 ] = 1'd1;
    assign memfont[655 ] = 1'd1;
    assign memfont[656 ] = 1'd1;
    assign memfont[657 ] = 1'd1;
    assign memfont[658 ] = 1'd1;
    assign memfont[659 ] = 1'd0;
    assign memfont[660 ] = 1'd0;
    assign memfont[661 ] = 1'd0;
    assign memfont[662 ] = 1'd0;
    assign memfont[663 ] = 1'd0;
    assign memfont[664 ] = 1'd0;
    assign memfont[665 ] = 1'd1;
    assign memfont[666 ] = 1'd1;
    assign memfont[667 ] = 1'd0;
    assign memfont[668 ] = 1'd0;
    assign memfont[669 ] = 1'd0;
    assign memfont[670 ] = 1'd0;
    assign memfont[671 ] = 1'd0;
    assign memfont[672 ] = 1'd0;
    assign memfont[673 ] = 1'd0;
    assign memfont[674 ] = 1'd0;
    assign memfont[675 ] = 1'd0;
    assign memfont[676 ] = 1'd0;
    assign memfont[677 ] = 1'd0;
    assign memfont[678 ] = 1'd0;
    assign memfont[679 ] = 1'd0;
    assign memfont[680 ] = 1'd0;
    assign memfont[681 ] = 1'd0;
    assign memfont[682 ] = 1'd0;
    assign memfont[683 ] = 1'd0;
    assign memfont[684 ] = 1'd0;
    assign memfont[685 ] = 1'd0;
    assign memfont[686 ] = 1'd0;
    assign memfont[687 ] = 1'd0;
    assign memfont[688 ] = 1'd0;
    assign memfont[689 ] = 1'd0;
    assign memfont[690 ] = 1'd0;
    assign memfont[691 ] = 1'd0;
    assign memfont[692 ] = 1'd0;
    assign memfont[693 ] = 1'd0;
    assign memfont[694 ] = 1'd0;
    assign memfont[695 ] = 1'd0;
    assign memfont[696 ] = 1'd0;
    assign memfont[697 ] = 1'd0;
    assign memfont[698 ] = 1'd0;
    assign memfont[699 ] = 1'd0;
    assign memfont[700 ] = 1'd0;
    assign memfont[701 ] = 1'd1;
    assign memfont[702 ] = 1'd1;
    assign memfont[703 ] = 1'd0;
    assign memfont[704 ] = 1'd0;
    assign memfont[705 ] = 1'd0;
    assign memfont[706 ] = 1'd0;
    assign memfont[707 ] = 1'd0;
    assign memfont[708 ] = 1'd0;
    assign memfont[709 ] = 1'd1;
    assign memfont[710 ] = 1'd1;
    assign memfont[711 ] = 1'd1;
    assign memfont[712 ] = 1'd1;
    assign memfont[713 ] = 1'd1;
    assign memfont[714 ] = 1'd1;
    assign memfont[715 ] = 1'd1;
    assign memfont[716 ] = 1'd1;
    assign memfont[717 ] = 1'd0;
    assign memfont[718 ] = 1'd0;
    assign memfont[719 ] = 1'd0;
    assign memfont[720 ] = 1'd0;
    assign memfont[721 ] = 1'd0;
    assign memfont[722 ] = 1'd0;
    assign memfont[723 ] = 1'd1;
    assign memfont[724 ] = 1'd1;
    assign memfont[725 ] = 1'd1;
    assign memfont[726 ] = 1'd1;
    assign memfont[727 ] = 1'd1;
    assign memfont[728 ] = 1'd1;
    assign memfont[729 ] = 1'd0;
    assign memfont[730 ] = 1'd0;
    assign memfont[731 ] = 1'd0;
    assign memfont[732 ] = 1'd0;
    assign memfont[733 ] = 1'd1;
    assign memfont[734 ] = 1'd1;
    assign memfont[735 ] = 1'd1;
    assign memfont[736 ] = 1'd1;
    assign memfont[737 ] = 1'd1;
    assign memfont[738 ] = 1'd1;
    assign memfont[739 ] = 1'd1;
    assign memfont[740 ] = 1'd0;
    assign memfont[741 ] = 1'd0;
    assign memfont[742 ] = 1'd0;
    assign memfont[743 ] = 1'd0;
    assign memfont[744 ] = 1'd0;
    assign memfont[745 ] = 1'd1;
    assign memfont[746 ] = 1'd1;
    assign memfont[747 ] = 1'd1;
    assign memfont[748 ] = 1'd1;
    assign memfont[749 ] = 1'd1;
    assign memfont[750 ] = 1'd1;
    assign memfont[751 ] = 1'd1;
    assign memfont[752 ] = 1'd1;
    assign memfont[753 ] = 1'd1;
    assign memfont[754 ] = 1'd0;
    assign memfont[755 ] = 1'd0;
    assign memfont[756 ] = 1'd0;
    assign memfont[757 ] = 1'd1;
    assign memfont[758 ] = 1'd1;
    assign memfont[759 ] = 1'd1;
    assign memfont[760 ] = 1'd1;
    assign memfont[761 ] = 1'd1;
    assign memfont[762 ] = 1'd1;
    assign memfont[763 ] = 1'd1;
    assign memfont[764 ] = 1'd1;
    assign memfont[765 ] = 1'd1;
    assign memfont[766 ] = 1'd1;
    assign memfont[767 ] = 1'd0;
    assign memfont[768 ] = 1'd0;
    assign memfont[769 ] = 1'd0;
    assign memfont[770 ] = 1'd0;
    assign memfont[771 ] = 1'd1;
    assign memfont[772 ] = 1'd1;
    assign memfont[773 ] = 1'd1;
    assign memfont[774 ] = 1'd1;
    assign memfont[775 ] = 1'd1;
    assign memfont[776 ] = 1'd1;
    assign memfont[777 ] = 1'd0;
    assign memfont[778 ] = 1'd0;
    assign memfont[779 ] = 1'd0;
    assign memfont[780 ] = 1'd0;
    assign memfont[781 ] = 1'd1;
    assign memfont[782 ] = 1'd1;
    assign memfont[783 ] = 1'd0;
    assign memfont[784 ] = 1'd0;
    assign memfont[785 ] = 1'd0;
    assign memfont[786 ] = 1'd0;
    assign memfont[787 ] = 1'd0;
    assign memfont[788 ] = 1'd0;
    assign memfont[789 ] = 1'd1;
    assign memfont[790 ] = 1'd1;
    assign memfont[791 ] = 1'd0;
    assign memfont[792 ] = 1'd0;
    assign memfont[793 ] = 1'd0;
    assign memfont[794 ] = 1'd0;
    assign memfont[795 ] = 1'd0;
    assign memfont[796 ] = 1'd0;
    assign memfont[797 ] = 1'd1;
    assign memfont[798 ] = 1'd1;
    assign memfont[799 ] = 1'd0;
    assign memfont[800 ] = 1'd0;
    assign memfont[801 ] = 1'd0;
    assign memfont[802 ] = 1'd0;
    assign memfont[803 ] = 1'd0;
    assign memfont[804 ] = 1'd0;
    assign memfont[805 ] = 1'd0;
    assign memfont[806 ] = 1'd0;
    assign memfont[807 ] = 1'd0;
    assign memfont[808 ] = 1'd0;
    assign memfont[809 ] = 1'd0;
    assign memfont[810 ] = 1'd0;
    assign memfont[811 ] = 1'd0;
    assign memfont[812 ] = 1'd1;
    assign memfont[813 ] = 1'd1;
    assign memfont[814 ] = 1'd1;
    assign memfont[815 ] = 1'd0;
    assign memfont[816 ] = 1'd0;
    assign memfont[817 ] = 1'd1;
    assign memfont[818 ] = 1'd1;
    assign memfont[819 ] = 1'd0;
    assign memfont[820 ] = 1'd0;
    assign memfont[821 ] = 1'd0;
    assign memfont[822 ] = 1'd0;
    assign memfont[823 ] = 1'd0;
    assign memfont[824 ] = 1'd1;
    assign memfont[825 ] = 1'd1;
    assign memfont[826 ] = 1'd0;
    assign memfont[827 ] = 1'd0;
    assign memfont[828 ] = 1'd0;
    assign memfont[829 ] = 1'd1;
    assign memfont[830 ] = 1'd1;
    assign memfont[831 ] = 1'd0;
    assign memfont[832 ] = 1'd0;
    assign memfont[833 ] = 1'd0;
    assign memfont[834 ] = 1'd0;
    assign memfont[835 ] = 1'd0;
    assign memfont[836 ] = 1'd0;
    assign memfont[837 ] = 1'd0;
    assign memfont[838 ] = 1'd0;
    assign memfont[839 ] = 1'd0;
    assign memfont[840 ] = 1'd0;
    assign memfont[841 ] = 1'd1;
    assign memfont[842 ] = 1'd1;
    assign memfont[843 ] = 1'd1;
    assign memfont[844 ] = 1'd0;
    assign memfont[845 ] = 1'd0;
    assign memfont[846 ] = 1'd0;
    assign memfont[847 ] = 1'd0;
    assign memfont[848 ] = 1'd1;
    assign memfont[849 ] = 1'd1;
    assign memfont[850 ] = 1'd1;
    assign memfont[851 ] = 1'd0;
    assign memfont[852 ] = 1'd0;
    assign memfont[853 ] = 1'd1;
    assign memfont[854 ] = 1'd1;
    assign memfont[855 ] = 1'd1;
    assign memfont[856 ] = 1'd0;
    assign memfont[857 ] = 1'd0;
    assign memfont[858 ] = 1'd0;
    assign memfont[859 ] = 1'd0;
    assign memfont[860 ] = 1'd0;
    assign memfont[861 ] = 1'd1;
    assign memfont[862 ] = 1'd1;
    assign memfont[863 ] = 1'd0;
    assign memfont[864 ] = 1'd0;
    assign memfont[865 ] = 1'd0;
    assign memfont[866 ] = 1'd0;
    assign memfont[867 ] = 1'd1;
    assign memfont[868 ] = 1'd1;
    assign memfont[869 ] = 1'd1;
    assign memfont[870 ] = 1'd1;
    assign memfont[871 ] = 1'd1;
    assign memfont[872 ] = 1'd1;
    assign memfont[873 ] = 1'd0;
    assign memfont[874 ] = 1'd0;
    assign memfont[875 ] = 1'd0;
    assign memfont[876 ] = 1'd0;
    assign memfont[877 ] = 1'd1;
    assign memfont[878 ] = 1'd1;
    assign memfont[879 ] = 1'd1;
    assign memfont[880 ] = 1'd1;
    assign memfont[881 ] = 1'd1;
    assign memfont[882 ] = 1'd1;
    assign memfont[883 ] = 1'd1;
    assign memfont[884 ] = 1'd1;
    assign memfont[885 ] = 1'd0;
    assign memfont[886 ] = 1'd0;
    assign memfont[887 ] = 1'd0;
    assign memfont[888 ] = 1'd0;
    assign memfont[889 ] = 1'd0;
    assign memfont[890 ] = 1'd0;
    assign memfont[891 ] = 1'd1;
    assign memfont[892 ] = 1'd1;
    assign memfont[893 ] = 1'd1;
    assign memfont[894 ] = 1'd1;
    assign memfont[895 ] = 1'd1;
    assign memfont[896 ] = 1'd1;
    assign memfont[897 ] = 1'd0;
    assign memfont[898 ] = 1'd0;
    assign memfont[899 ] = 1'd0;
    assign memfont[900 ] = 1'd0;
    assign memfont[901 ] = 1'd1;
    assign memfont[902 ] = 1'd1;
    assign memfont[903 ] = 1'd1;
    assign memfont[904 ] = 1'd1;
    assign memfont[905 ] = 1'd1;
    assign memfont[906 ] = 1'd1;
    assign memfont[907 ] = 1'd1;
    assign memfont[908 ] = 1'd1;
    assign memfont[909 ] = 1'd0;
    assign memfont[910 ] = 1'd0;
    assign memfont[911 ] = 1'd0;
    assign memfont[912 ] = 1'd0;
    assign memfont[913 ] = 1'd0;
    assign memfont[914 ] = 1'd0;
    assign memfont[915 ] = 1'd1;
    assign memfont[916 ] = 1'd1;
    assign memfont[917 ] = 1'd1;
    assign memfont[918 ] = 1'd1;
    assign memfont[919 ] = 1'd1;
    assign memfont[920 ] = 1'd1;
    assign memfont[921 ] = 1'd0;
    assign memfont[922 ] = 1'd0;
    assign memfont[923 ] = 1'd0;
    assign memfont[924 ] = 1'd0;
    assign memfont[925 ] = 1'd1;
    assign memfont[926 ] = 1'd1;
    assign memfont[927 ] = 1'd1;
    assign memfont[928 ] = 1'd1;
    assign memfont[929 ] = 1'd1;
    assign memfont[930 ] = 1'd1;
    assign memfont[931 ] = 1'd1;
    assign memfont[932 ] = 1'd1;
    assign memfont[933 ] = 1'd1;
    assign memfont[934 ] = 1'd1;
    assign memfont[935 ] = 1'd0;
    assign memfont[936 ] = 1'd0;
    assign memfont[937 ] = 1'd1;
    assign memfont[938 ] = 1'd1;
    assign memfont[939 ] = 1'd0;
    assign memfont[940 ] = 1'd0;
    assign memfont[941 ] = 1'd0;
    assign memfont[942 ] = 1'd0;
    assign memfont[943 ] = 1'd0;
    assign memfont[944 ] = 1'd0;
    assign memfont[945 ] = 1'd1;
    assign memfont[946 ] = 1'd1;
    assign memfont[947 ] = 1'd0;
    assign memfont[948 ] = 1'd1;
    assign memfont[949 ] = 1'd1;
    assign memfont[950 ] = 1'd1;
    assign memfont[951 ] = 1'd0;
    assign memfont[952 ] = 1'd0;
    assign memfont[953 ] = 1'd0;
    assign memfont[954 ] = 1'd0;
    assign memfont[955 ] = 1'd0;
    assign memfont[956 ] = 1'd0;
    assign memfont[957 ] = 1'd1;
    assign memfont[958 ] = 1'd1;
    assign memfont[959 ] = 1'd0;
    assign memfont[960 ] = 1'd1;
    assign memfont[961 ] = 1'd1;
    assign memfont[962 ] = 1'd0;
    assign memfont[963 ] = 1'd0;
    assign memfont[964 ] = 1'd0;
    assign memfont[965 ] = 1'd1;
    assign memfont[966 ] = 1'd1;
    assign memfont[967 ] = 1'd0;
    assign memfont[968 ] = 1'd0;
    assign memfont[969 ] = 1'd1;
    assign memfont[970 ] = 1'd1;
    assign memfont[971 ] = 1'd0;
    assign memfont[972 ] = 1'd0;
    assign memfont[973 ] = 1'd1;
    assign memfont[974 ] = 1'd1;
    assign memfont[975 ] = 1'd1;
    assign memfont[976 ] = 1'd0;
    assign memfont[977 ] = 1'd0;
    assign memfont[978 ] = 1'd0;
    assign memfont[979 ] = 1'd0;
    assign memfont[980 ] = 1'd1;
    assign memfont[981 ] = 1'd1;
    assign memfont[982 ] = 1'd0;
    assign memfont[983 ] = 1'd0;
    assign memfont[984 ] = 1'd0;
    assign memfont[985 ] = 1'd1;
    assign memfont[986 ] = 1'd1;
    assign memfont[987 ] = 1'd0;
    assign memfont[988 ] = 1'd0;
    assign memfont[989 ] = 1'd0;
    assign memfont[990 ] = 1'd0;
    assign memfont[991 ] = 1'd0;
    assign memfont[992 ] = 1'd0;
    assign memfont[993 ] = 1'd1;
    assign memfont[994 ] = 1'd1;
    assign memfont[995 ] = 1'd0;
    assign memfont[996 ] = 1'd0;
    assign memfont[997 ] = 1'd1;
    assign memfont[998 ] = 1'd1;
    assign memfont[999 ] = 1'd1;
    assign memfont[1000] = 1'd1;
    assign memfont[1001] = 1'd1;
    assign memfont[1002] = 1'd1;
    assign memfont[1003] = 1'd1;
    assign memfont[1004] = 1'd1;
    assign memfont[1005] = 1'd1;
    assign memfont[1006] = 1'd1;
    assign memfont[1007] = 1'd0;
    assign memfont[1008] = 1'd0;
    assign memfont[1009] = 1'd0;
    assign memfont[1010] = 1'd0;
    assign memfont[1011] = 1'd0;
    assign memfont[1012] = 1'd0;
    assign memfont[1013] = 1'd1;
    assign memfont[1014] = 1'd1;
    assign memfont[1015] = 1'd0;
    assign memfont[1016] = 1'd0;
    assign memfont[1017] = 1'd0;
    assign memfont[1018] = 1'd0;
    assign memfont[1019] = 1'd0;
    assign memfont[1020] = 1'd0;
    assign memfont[1021] = 1'd0;
    assign memfont[1022] = 1'd0;
    assign memfont[1023] = 1'd0;
    assign memfont[1024] = 1'd0;
    assign memfont[1025] = 1'd0;
    assign memfont[1026] = 1'd0;
    assign memfont[1027] = 1'd0;
    assign memfont[1028] = 1'd0;
    assign memfont[1029] = 1'd0;
    assign memfont[1030] = 1'd0;
    assign memfont[1031] = 1'd0;
    assign memfont[1032] = 1'd0;
    assign memfont[1033] = 1'd0;
    assign memfont[1034] = 1'd0;
    assign memfont[1035] = 1'd0;
    assign memfont[1036] = 1'd0;
    assign memfont[1037] = 1'd0;
    assign memfont[1038] = 1'd0;
    assign memfont[1039] = 1'd0;
    assign memfont[1040] = 1'd0;
    assign memfont[1041] = 1'd0;
    assign memfont[1042] = 1'd0;
    assign memfont[1043] = 1'd0;
    assign memfont[1044] = 1'd0;
    assign memfont[1045] = 1'd0;
    assign memfont[1046] = 1'd0;
    assign memfont[1047] = 1'd0;
    assign memfont[1048] = 1'd1;
    assign memfont[1049] = 1'd1;
    assign memfont[1050] = 1'd1;
    assign memfont[1051] = 1'd0;
    assign memfont[1052] = 1'd0;
    assign memfont[1053] = 1'd0;
    assign memfont[1054] = 1'd0;
    assign memfont[1055] = 1'd0;
    assign memfont[1056] = 1'd0;
    assign memfont[1057] = 1'd1;
    assign memfont[1058] = 1'd1;
    assign memfont[1059] = 1'd0;
    assign memfont[1060] = 1'd0;
    assign memfont[1061] = 1'd0;
    assign memfont[1062] = 1'd0;
    assign memfont[1063] = 1'd1;
    assign memfont[1064] = 1'd1;
    assign memfont[1065] = 1'd1;
    assign memfont[1066] = 1'd0;
    assign memfont[1067] = 1'd0;
    assign memfont[1068] = 1'd0;
    assign memfont[1069] = 1'd0;
    assign memfont[1070] = 1'd1;
    assign memfont[1071] = 1'd1;
    assign memfont[1072] = 1'd1;
    assign memfont[1073] = 1'd0;
    assign memfont[1074] = 1'd0;
    assign memfont[1075] = 1'd0;
    assign memfont[1076] = 1'd1;
    assign memfont[1077] = 1'd1;
    assign memfont[1078] = 1'd0;
    assign memfont[1079] = 1'd0;
    assign memfont[1080] = 1'd0;
    assign memfont[1081] = 1'd1;
    assign memfont[1082] = 1'd1;
    assign memfont[1083] = 1'd0;
    assign memfont[1084] = 1'd0;
    assign memfont[1085] = 1'd0;
    assign memfont[1086] = 1'd1;
    assign memfont[1087] = 1'd1;
    assign memfont[1088] = 1'd1;
    assign memfont[1089] = 1'd0;
    assign memfont[1090] = 1'd0;
    assign memfont[1091] = 1'd0;
    assign memfont[1092] = 1'd0;
    assign memfont[1093] = 1'd1;
    assign memfont[1094] = 1'd1;
    assign memfont[1095] = 1'd0;
    assign memfont[1096] = 1'd0;
    assign memfont[1097] = 1'd0;
    assign memfont[1098] = 1'd0;
    assign memfont[1099] = 1'd0;
    assign memfont[1100] = 1'd0;
    assign memfont[1101] = 1'd0;
    assign memfont[1102] = 1'd0;
    assign memfont[1103] = 1'd0;
    assign memfont[1104] = 1'd0;
    assign memfont[1105] = 1'd1;
    assign memfont[1106] = 1'd1;
    assign memfont[1107] = 1'd0;
    assign memfont[1108] = 1'd0;
    assign memfont[1109] = 1'd0;
    assign memfont[1110] = 1'd0;
    assign memfont[1111] = 1'd0;
    assign memfont[1112] = 1'd0;
    assign memfont[1113] = 1'd0;
    assign memfont[1114] = 1'd0;
    assign memfont[1115] = 1'd0;
    assign memfont[1116] = 1'd0;
    assign memfont[1117] = 1'd0;
    assign memfont[1118] = 1'd1;
    assign memfont[1119] = 1'd1;
    assign memfont[1120] = 1'd1;
    assign memfont[1121] = 1'd0;
    assign memfont[1122] = 1'd0;
    assign memfont[1123] = 1'd1;
    assign memfont[1124] = 1'd1;
    assign memfont[1125] = 1'd1;
    assign memfont[1126] = 1'd0;
    assign memfont[1127] = 1'd0;
    assign memfont[1128] = 1'd0;
    assign memfont[1129] = 1'd1;
    assign memfont[1130] = 1'd1;
    assign memfont[1131] = 1'd0;
    assign memfont[1132] = 1'd0;
    assign memfont[1133] = 1'd0;
    assign memfont[1134] = 1'd0;
    assign memfont[1135] = 1'd0;
    assign memfont[1136] = 1'd0;
    assign memfont[1137] = 1'd1;
    assign memfont[1138] = 1'd1;
    assign memfont[1139] = 1'd0;
    assign memfont[1140] = 1'd0;
    assign memfont[1141] = 1'd0;
    assign memfont[1142] = 1'd0;
    assign memfont[1143] = 1'd0;
    assign memfont[1144] = 1'd0;
    assign memfont[1145] = 1'd1;
    assign memfont[1146] = 1'd1;
    assign memfont[1147] = 1'd0;
    assign memfont[1148] = 1'd0;
    assign memfont[1149] = 1'd0;
    assign memfont[1150] = 1'd0;
    assign memfont[1151] = 1'd0;
    assign memfont[1152] = 1'd0;
    assign memfont[1153] = 1'd0;
    assign memfont[1154] = 1'd0;
    assign memfont[1155] = 1'd0;
    assign memfont[1156] = 1'd0;
    assign memfont[1157] = 1'd0;
    assign memfont[1158] = 1'd0;
    assign memfont[1159] = 1'd0;
    assign memfont[1160] = 1'd1;
    assign memfont[1161] = 1'd1;
    assign memfont[1162] = 1'd1;
    assign memfont[1163] = 1'd0;
    assign memfont[1164] = 1'd0;
    assign memfont[1165] = 1'd1;
    assign memfont[1166] = 1'd1;
    assign memfont[1167] = 1'd0;
    assign memfont[1168] = 1'd0;
    assign memfont[1169] = 1'd0;
    assign memfont[1170] = 1'd0;
    assign memfont[1171] = 1'd1;
    assign memfont[1172] = 1'd1;
    assign memfont[1173] = 1'd0;
    assign memfont[1174] = 1'd0;
    assign memfont[1175] = 1'd0;
    assign memfont[1176] = 1'd0;
    assign memfont[1177] = 1'd1;
    assign memfont[1178] = 1'd1;
    assign memfont[1179] = 1'd0;
    assign memfont[1180] = 1'd0;
    assign memfont[1181] = 1'd0;
    assign memfont[1182] = 1'd0;
    assign memfont[1183] = 1'd0;
    assign memfont[1184] = 1'd0;
    assign memfont[1185] = 1'd0;
    assign memfont[1186] = 1'd0;
    assign memfont[1187] = 1'd0;
    assign memfont[1188] = 1'd0;
    assign memfont[1189] = 1'd1;
    assign memfont[1190] = 1'd1;
    assign memfont[1191] = 1'd1;
    assign memfont[1192] = 1'd0;
    assign memfont[1193] = 1'd0;
    assign memfont[1194] = 1'd0;
    assign memfont[1195] = 1'd0;
    assign memfont[1196] = 1'd1;
    assign memfont[1197] = 1'd1;
    assign memfont[1198] = 1'd1;
    assign memfont[1199] = 1'd0;
    assign memfont[1200] = 1'd0;
    assign memfont[1201] = 1'd1;
    assign memfont[1202] = 1'd1;
    assign memfont[1203] = 1'd1;
    assign memfont[1204] = 1'd0;
    assign memfont[1205] = 1'd0;
    assign memfont[1206] = 1'd0;
    assign memfont[1207] = 1'd0;
    assign memfont[1208] = 1'd0;
    assign memfont[1209] = 1'd1;
    assign memfont[1210] = 1'd1;
    assign memfont[1211] = 1'd0;
    assign memfont[1212] = 1'd0;
    assign memfont[1213] = 1'd0;
    assign memfont[1214] = 1'd1;
    assign memfont[1215] = 1'd1;
    assign memfont[1216] = 1'd1;
    assign memfont[1217] = 1'd0;
    assign memfont[1218] = 1'd0;
    assign memfont[1219] = 1'd1;
    assign memfont[1220] = 1'd1;
    assign memfont[1221] = 1'd1;
    assign memfont[1222] = 1'd0;
    assign memfont[1223] = 1'd0;
    assign memfont[1224] = 1'd0;
    assign memfont[1225] = 1'd1;
    assign memfont[1226] = 1'd1;
    assign memfont[1227] = 1'd0;
    assign memfont[1228] = 1'd0;
    assign memfont[1229] = 1'd0;
    assign memfont[1230] = 1'd0;
    assign memfont[1231] = 1'd1;
    assign memfont[1232] = 1'd1;
    assign memfont[1233] = 1'd1;
    assign memfont[1234] = 1'd0;
    assign memfont[1235] = 1'd0;
    assign memfont[1236] = 1'd0;
    assign memfont[1237] = 1'd0;
    assign memfont[1238] = 1'd1;
    assign memfont[1239] = 1'd1;
    assign memfont[1240] = 1'd1;
    assign memfont[1241] = 1'd0;
    assign memfont[1242] = 1'd0;
    assign memfont[1243] = 1'd1;
    assign memfont[1244] = 1'd1;
    assign memfont[1245] = 1'd1;
    assign memfont[1246] = 1'd0;
    assign memfont[1247] = 1'd0;
    assign memfont[1248] = 1'd0;
    assign memfont[1249] = 1'd1;
    assign memfont[1250] = 1'd1;
    assign memfont[1251] = 1'd0;
    assign memfont[1252] = 1'd0;
    assign memfont[1253] = 1'd0;
    assign memfont[1254] = 1'd0;
    assign memfont[1255] = 1'd1;
    assign memfont[1256] = 1'd1;
    assign memfont[1257] = 1'd1;
    assign memfont[1258] = 1'd0;
    assign memfont[1259] = 1'd0;
    assign memfont[1260] = 1'd0;
    assign memfont[1261] = 1'd0;
    assign memfont[1262] = 1'd1;
    assign memfont[1263] = 1'd1;
    assign memfont[1264] = 1'd0;
    assign memfont[1265] = 1'd0;
    assign memfont[1266] = 1'd0;
    assign memfont[1267] = 1'd1;
    assign memfont[1268] = 1'd1;
    assign memfont[1269] = 1'd1;
    assign memfont[1270] = 1'd0;
    assign memfont[1271] = 1'd0;
    assign memfont[1272] = 1'd0;
    assign memfont[1273] = 1'd0;
    assign memfont[1274] = 1'd0;
    assign memfont[1275] = 1'd0;
    assign memfont[1276] = 1'd0;
    assign memfont[1277] = 1'd1;
    assign memfont[1278] = 1'd1;
    assign memfont[1279] = 1'd0;
    assign memfont[1280] = 1'd0;
    assign memfont[1281] = 1'd0;
    assign memfont[1282] = 1'd0;
    assign memfont[1283] = 1'd0;
    assign memfont[1284] = 1'd0;
    assign memfont[1285] = 1'd1;
    assign memfont[1286] = 1'd1;
    assign memfont[1287] = 1'd0;
    assign memfont[1288] = 1'd0;
    assign memfont[1289] = 1'd0;
    assign memfont[1290] = 1'd0;
    assign memfont[1291] = 1'd0;
    assign memfont[1292] = 1'd0;
    assign memfont[1293] = 1'd1;
    assign memfont[1294] = 1'd1;
    assign memfont[1295] = 1'd0;
    assign memfont[1296] = 1'd0;
    assign memfont[1297] = 1'd1;
    assign memfont[1298] = 1'd1;
    assign memfont[1299] = 1'd0;
    assign memfont[1300] = 1'd0;
    assign memfont[1301] = 1'd0;
    assign memfont[1302] = 1'd0;
    assign memfont[1303] = 1'd0;
    assign memfont[1304] = 1'd0;
    assign memfont[1305] = 1'd1;
    assign memfont[1306] = 1'd1;
    assign memfont[1307] = 1'd0;
    assign memfont[1308] = 1'd1;
    assign memfont[1309] = 1'd1;
    assign memfont[1310] = 1'd0;
    assign memfont[1311] = 1'd0;
    assign memfont[1312] = 1'd0;
    assign memfont[1313] = 1'd1;
    assign memfont[1314] = 1'd1;
    assign memfont[1315] = 1'd0;
    assign memfont[1316] = 1'd0;
    assign memfont[1317] = 1'd1;
    assign memfont[1318] = 1'd1;
    assign memfont[1319] = 1'd0;
    assign memfont[1320] = 1'd0;
    assign memfont[1321] = 1'd0;
    assign memfont[1322] = 1'd1;
    assign memfont[1323] = 1'd1;
    assign memfont[1324] = 1'd0;
    assign memfont[1325] = 1'd0;
    assign memfont[1326] = 1'd0;
    assign memfont[1327] = 1'd0;
    assign memfont[1328] = 1'd1;
    assign memfont[1329] = 1'd1;
    assign memfont[1330] = 1'd0;
    assign memfont[1331] = 1'd0;
    assign memfont[1332] = 1'd0;
    assign memfont[1333] = 1'd1;
    assign memfont[1334] = 1'd1;
    assign memfont[1335] = 1'd0;
    assign memfont[1336] = 1'd0;
    assign memfont[1337] = 1'd0;
    assign memfont[1338] = 1'd0;
    assign memfont[1339] = 1'd0;
    assign memfont[1340] = 1'd1;
    assign memfont[1341] = 1'd1;
    assign memfont[1342] = 1'd0;
    assign memfont[1343] = 1'd0;
    assign memfont[1344] = 1'd0;
    assign memfont[1345] = 1'd0;
    assign memfont[1346] = 1'd0;
    assign memfont[1347] = 1'd0;
    assign memfont[1348] = 1'd0;
    assign memfont[1349] = 1'd0;
    assign memfont[1350] = 1'd0;
    assign memfont[1351] = 1'd0;
    assign memfont[1352] = 1'd1;
    assign memfont[1353] = 1'd1;
    assign memfont[1354] = 1'd0;
    assign memfont[1355] = 1'd0;
    assign memfont[1356] = 1'd0;
    assign memfont[1357] = 1'd0;
    assign memfont[1358] = 1'd0;
    assign memfont[1359] = 1'd0;
    assign memfont[1360] = 1'd0;
    assign memfont[1361] = 1'd1;
    assign memfont[1362] = 1'd1;
    assign memfont[1363] = 1'd0;
    assign memfont[1364] = 1'd0;
    assign memfont[1365] = 1'd0;
    assign memfont[1366] = 1'd0;
    assign memfont[1367] = 1'd0;
    assign memfont[1368] = 1'd0;
    assign memfont[1369] = 1'd0;
    assign memfont[1370] = 1'd0;
    assign memfont[1371] = 1'd0;
    assign memfont[1372] = 1'd0;
    assign memfont[1373] = 1'd0;
    assign memfont[1374] = 1'd0;
    assign memfont[1375] = 1'd0;
    assign memfont[1376] = 1'd0;
    assign memfont[1377] = 1'd0;
    assign memfont[1378] = 1'd0;
    assign memfont[1379] = 1'd0;
    assign memfont[1380] = 1'd0;
    assign memfont[1381] = 1'd0;
    assign memfont[1382] = 1'd0;
    assign memfont[1383] = 1'd0;
    assign memfont[1384] = 1'd0;
    assign memfont[1385] = 1'd0;
    assign memfont[1386] = 1'd0;
    assign memfont[1387] = 1'd0;
    assign memfont[1388] = 1'd0;
    assign memfont[1389] = 1'd0;
    assign memfont[1390] = 1'd0;
    assign memfont[1391] = 1'd0;
    assign memfont[1392] = 1'd0;
    assign memfont[1393] = 1'd0;
    assign memfont[1394] = 1'd0;
    assign memfont[1395] = 1'd0;
    assign memfont[1396] = 1'd1;
    assign memfont[1397] = 1'd1;
    assign memfont[1398] = 1'd1;
    assign memfont[1399] = 1'd1;
    assign memfont[1400] = 1'd0;
    assign memfont[1401] = 1'd0;
    assign memfont[1402] = 1'd0;
    assign memfont[1403] = 1'd0;
    assign memfont[1404] = 1'd0;
    assign memfont[1405] = 1'd1;
    assign memfont[1406] = 1'd1;
    assign memfont[1407] = 1'd0;
    assign memfont[1408] = 1'd0;
    assign memfont[1409] = 1'd0;
    assign memfont[1410] = 1'd0;
    assign memfont[1411] = 1'd0;
    assign memfont[1412] = 1'd1;
    assign memfont[1413] = 1'd1;
    assign memfont[1414] = 1'd0;
    assign memfont[1415] = 1'd0;
    assign memfont[1416] = 1'd0;
    assign memfont[1417] = 1'd0;
    assign memfont[1418] = 1'd1;
    assign memfont[1419] = 1'd1;
    assign memfont[1420] = 1'd0;
    assign memfont[1421] = 1'd0;
    assign memfont[1422] = 1'd0;
    assign memfont[1423] = 1'd0;
    assign memfont[1424] = 1'd0;
    assign memfont[1425] = 1'd1;
    assign memfont[1426] = 1'd1;
    assign memfont[1427] = 1'd0;
    assign memfont[1428] = 1'd0;
    assign memfont[1429] = 1'd1;
    assign memfont[1430] = 1'd1;
    assign memfont[1431] = 1'd0;
    assign memfont[1432] = 1'd0;
    assign memfont[1433] = 1'd0;
    assign memfont[1434] = 1'd0;
    assign memfont[1435] = 1'd1;
    assign memfont[1436] = 1'd1;
    assign memfont[1437] = 1'd1;
    assign memfont[1438] = 1'd0;
    assign memfont[1439] = 1'd0;
    assign memfont[1440] = 1'd0;
    assign memfont[1441] = 1'd1;
    assign memfont[1442] = 1'd1;
    assign memfont[1443] = 1'd0;
    assign memfont[1444] = 1'd0;
    assign memfont[1445] = 1'd0;
    assign memfont[1446] = 1'd0;
    assign memfont[1447] = 1'd0;
    assign memfont[1448] = 1'd0;
    assign memfont[1449] = 1'd0;
    assign memfont[1450] = 1'd0;
    assign memfont[1451] = 1'd0;
    assign memfont[1452] = 1'd0;
    assign memfont[1453] = 1'd1;
    assign memfont[1454] = 1'd1;
    assign memfont[1455] = 1'd0;
    assign memfont[1456] = 1'd0;
    assign memfont[1457] = 1'd0;
    assign memfont[1458] = 1'd0;
    assign memfont[1459] = 1'd0;
    assign memfont[1460] = 1'd0;
    assign memfont[1461] = 1'd0;
    assign memfont[1462] = 1'd0;
    assign memfont[1463] = 1'd0;
    assign memfont[1464] = 1'd0;
    assign memfont[1465] = 1'd0;
    assign memfont[1466] = 1'd1;
    assign memfont[1467] = 1'd1;
    assign memfont[1468] = 1'd0;
    assign memfont[1469] = 1'd0;
    assign memfont[1470] = 1'd0;
    assign memfont[1471] = 1'd0;
    assign memfont[1472] = 1'd1;
    assign memfont[1473] = 1'd1;
    assign memfont[1474] = 1'd0;
    assign memfont[1475] = 1'd0;
    assign memfont[1476] = 1'd0;
    assign memfont[1477] = 1'd1;
    assign memfont[1478] = 1'd1;
    assign memfont[1479] = 1'd0;
    assign memfont[1480] = 1'd0;
    assign memfont[1481] = 1'd0;
    assign memfont[1482] = 1'd0;
    assign memfont[1483] = 1'd0;
    assign memfont[1484] = 1'd0;
    assign memfont[1485] = 1'd1;
    assign memfont[1486] = 1'd1;
    assign memfont[1487] = 1'd0;
    assign memfont[1488] = 1'd0;
    assign memfont[1489] = 1'd0;
    assign memfont[1490] = 1'd0;
    assign memfont[1491] = 1'd0;
    assign memfont[1492] = 1'd0;
    assign memfont[1493] = 1'd1;
    assign memfont[1494] = 1'd1;
    assign memfont[1495] = 1'd0;
    assign memfont[1496] = 1'd0;
    assign memfont[1497] = 1'd0;
    assign memfont[1498] = 1'd0;
    assign memfont[1499] = 1'd0;
    assign memfont[1500] = 1'd0;
    assign memfont[1501] = 1'd0;
    assign memfont[1502] = 1'd0;
    assign memfont[1503] = 1'd0;
    assign memfont[1504] = 1'd0;
    assign memfont[1505] = 1'd0;
    assign memfont[1506] = 1'd0;
    assign memfont[1507] = 1'd0;
    assign memfont[1508] = 1'd1;
    assign memfont[1509] = 1'd1;
    assign memfont[1510] = 1'd1;
    assign memfont[1511] = 1'd0;
    assign memfont[1512] = 1'd0;
    assign memfont[1513] = 1'd1;
    assign memfont[1514] = 1'd1;
    assign memfont[1515] = 1'd0;
    assign memfont[1516] = 1'd0;
    assign memfont[1517] = 1'd0;
    assign memfont[1518] = 1'd1;
    assign memfont[1519] = 1'd1;
    assign memfont[1520] = 1'd1;
    assign memfont[1521] = 1'd0;
    assign memfont[1522] = 1'd0;
    assign memfont[1523] = 1'd0;
    assign memfont[1524] = 1'd0;
    assign memfont[1525] = 1'd1;
    assign memfont[1526] = 1'd1;
    assign memfont[1527] = 1'd0;
    assign memfont[1528] = 1'd0;
    assign memfont[1529] = 1'd0;
    assign memfont[1530] = 1'd0;
    assign memfont[1531] = 1'd0;
    assign memfont[1532] = 1'd0;
    assign memfont[1533] = 1'd0;
    assign memfont[1534] = 1'd0;
    assign memfont[1535] = 1'd0;
    assign memfont[1536] = 1'd0;
    assign memfont[1537] = 1'd1;
    assign memfont[1538] = 1'd1;
    assign memfont[1539] = 1'd1;
    assign memfont[1540] = 1'd0;
    assign memfont[1541] = 1'd0;
    assign memfont[1542] = 1'd0;
    assign memfont[1543] = 1'd1;
    assign memfont[1544] = 1'd1;
    assign memfont[1545] = 1'd1;
    assign memfont[1546] = 1'd1;
    assign memfont[1547] = 1'd0;
    assign memfont[1548] = 1'd0;
    assign memfont[1549] = 1'd1;
    assign memfont[1550] = 1'd1;
    assign memfont[1551] = 1'd1;
    assign memfont[1552] = 1'd1;
    assign memfont[1553] = 1'd0;
    assign memfont[1554] = 1'd0;
    assign memfont[1555] = 1'd0;
    assign memfont[1556] = 1'd0;
    assign memfont[1557] = 1'd1;
    assign memfont[1558] = 1'd1;
    assign memfont[1559] = 1'd0;
    assign memfont[1560] = 1'd0;
    assign memfont[1561] = 1'd1;
    assign memfont[1562] = 1'd1;
    assign memfont[1563] = 1'd1;
    assign memfont[1564] = 1'd0;
    assign memfont[1565] = 1'd0;
    assign memfont[1566] = 1'd0;
    assign memfont[1567] = 1'd0;
    assign memfont[1568] = 1'd1;
    assign memfont[1569] = 1'd1;
    assign memfont[1570] = 1'd0;
    assign memfont[1571] = 1'd0;
    assign memfont[1572] = 1'd0;
    assign memfont[1573] = 1'd1;
    assign memfont[1574] = 1'd1;
    assign memfont[1575] = 1'd0;
    assign memfont[1576] = 1'd0;
    assign memfont[1577] = 1'd0;
    assign memfont[1578] = 1'd0;
    assign memfont[1579] = 1'd0;
    assign memfont[1580] = 1'd0;
    assign memfont[1581] = 1'd1;
    assign memfont[1582] = 1'd1;
    assign memfont[1583] = 1'd0;
    assign memfont[1584] = 1'd0;
    assign memfont[1585] = 1'd1;
    assign memfont[1586] = 1'd1;
    assign memfont[1587] = 1'd1;
    assign memfont[1588] = 1'd0;
    assign memfont[1589] = 1'd0;
    assign memfont[1590] = 1'd0;
    assign memfont[1591] = 1'd0;
    assign memfont[1592] = 1'd1;
    assign memfont[1593] = 1'd1;
    assign memfont[1594] = 1'd0;
    assign memfont[1595] = 1'd0;
    assign memfont[1596] = 1'd0;
    assign memfont[1597] = 1'd1;
    assign memfont[1598] = 1'd1;
    assign memfont[1599] = 1'd0;
    assign memfont[1600] = 1'd0;
    assign memfont[1601] = 1'd0;
    assign memfont[1602] = 1'd0;
    assign memfont[1603] = 1'd0;
    assign memfont[1604] = 1'd1;
    assign memfont[1605] = 1'd1;
    assign memfont[1606] = 1'd1;
    assign memfont[1607] = 1'd0;
    assign memfont[1608] = 1'd0;
    assign memfont[1609] = 1'd1;
    assign memfont[1610] = 1'd1;
    assign memfont[1611] = 1'd1;
    assign memfont[1612] = 1'd0;
    assign memfont[1613] = 1'd0;
    assign memfont[1614] = 1'd0;
    assign memfont[1615] = 1'd0;
    assign memfont[1616] = 1'd1;
    assign memfont[1617] = 1'd1;
    assign memfont[1618] = 1'd0;
    assign memfont[1619] = 1'd0;
    assign memfont[1620] = 1'd0;
    assign memfont[1621] = 1'd0;
    assign memfont[1622] = 1'd0;
    assign memfont[1623] = 1'd0;
    assign memfont[1624] = 1'd0;
    assign memfont[1625] = 1'd1;
    assign memfont[1626] = 1'd1;
    assign memfont[1627] = 1'd0;
    assign memfont[1628] = 1'd0;
    assign memfont[1629] = 1'd0;
    assign memfont[1630] = 1'd0;
    assign memfont[1631] = 1'd0;
    assign memfont[1632] = 1'd0;
    assign memfont[1633] = 1'd1;
    assign memfont[1634] = 1'd1;
    assign memfont[1635] = 1'd0;
    assign memfont[1636] = 1'd0;
    assign memfont[1637] = 1'd0;
    assign memfont[1638] = 1'd0;
    assign memfont[1639] = 1'd0;
    assign memfont[1640] = 1'd0;
    assign memfont[1641] = 1'd1;
    assign memfont[1642] = 1'd1;
    assign memfont[1643] = 1'd0;
    assign memfont[1644] = 1'd0;
    assign memfont[1645] = 1'd1;
    assign memfont[1646] = 1'd1;
    assign memfont[1647] = 1'd0;
    assign memfont[1648] = 1'd0;
    assign memfont[1649] = 1'd0;
    assign memfont[1650] = 1'd0;
    assign memfont[1651] = 1'd0;
    assign memfont[1652] = 1'd1;
    assign memfont[1653] = 1'd1;
    assign memfont[1654] = 1'd1;
    assign memfont[1655] = 1'd0;
    assign memfont[1656] = 1'd1;
    assign memfont[1657] = 1'd1;
    assign memfont[1658] = 1'd0;
    assign memfont[1659] = 1'd0;
    assign memfont[1660] = 1'd1;
    assign memfont[1661] = 1'd1;
    assign memfont[1662] = 1'd1;
    assign memfont[1663] = 1'd0;
    assign memfont[1664] = 1'd0;
    assign memfont[1665] = 1'd1;
    assign memfont[1666] = 1'd1;
    assign memfont[1667] = 1'd0;
    assign memfont[1668] = 1'd0;
    assign memfont[1669] = 1'd0;
    assign memfont[1670] = 1'd1;
    assign memfont[1671] = 1'd1;
    assign memfont[1672] = 1'd0;
    assign memfont[1673] = 1'd0;
    assign memfont[1674] = 1'd0;
    assign memfont[1675] = 1'd1;
    assign memfont[1676] = 1'd1;
    assign memfont[1677] = 1'd0;
    assign memfont[1678] = 1'd0;
    assign memfont[1679] = 1'd0;
    assign memfont[1680] = 1'd0;
    assign memfont[1681] = 1'd0;
    assign memfont[1682] = 1'd1;
    assign memfont[1683] = 1'd1;
    assign memfont[1684] = 1'd0;
    assign memfont[1685] = 1'd0;
    assign memfont[1686] = 1'd0;
    assign memfont[1687] = 1'd0;
    assign memfont[1688] = 1'd1;
    assign memfont[1689] = 1'd1;
    assign memfont[1690] = 1'd0;
    assign memfont[1691] = 1'd0;
    assign memfont[1692] = 1'd0;
    assign memfont[1693] = 1'd0;
    assign memfont[1694] = 1'd0;
    assign memfont[1695] = 1'd0;
    assign memfont[1696] = 1'd0;
    assign memfont[1697] = 1'd0;
    assign memfont[1698] = 1'd0;
    assign memfont[1699] = 1'd0;
    assign memfont[1700] = 1'd1;
    assign memfont[1701] = 1'd1;
    assign memfont[1702] = 1'd0;
    assign memfont[1703] = 1'd0;
    assign memfont[1704] = 1'd0;
    assign memfont[1705] = 1'd0;
    assign memfont[1706] = 1'd0;
    assign memfont[1707] = 1'd0;
    assign memfont[1708] = 1'd0;
    assign memfont[1709] = 1'd1;
    assign memfont[1710] = 1'd1;
    assign memfont[1711] = 1'd0;
    assign memfont[1712] = 1'd0;
    assign memfont[1713] = 1'd0;
    assign memfont[1714] = 1'd0;
    assign memfont[1715] = 1'd0;
    assign memfont[1716] = 1'd0;
    assign memfont[1717] = 1'd1;
    assign memfont[1718] = 1'd1;
    assign memfont[1719] = 1'd1;
    assign memfont[1720] = 1'd1;
    assign memfont[1721] = 1'd1;
    assign memfont[1722] = 1'd1;
    assign memfont[1723] = 1'd1;
    assign memfont[1724] = 1'd1;
    assign memfont[1725] = 1'd1;
    assign memfont[1726] = 1'd1;
    assign memfont[1727] = 1'd0;
    assign memfont[1728] = 1'd0;
    assign memfont[1729] = 1'd1;
    assign memfont[1730] = 1'd1;
    assign memfont[1731] = 1'd1;
    assign memfont[1732] = 1'd1;
    assign memfont[1733] = 1'd1;
    assign memfont[1734] = 1'd1;
    assign memfont[1735] = 1'd1;
    assign memfont[1736] = 1'd1;
    assign memfont[1737] = 1'd1;
    assign memfont[1738] = 1'd1;
    assign memfont[1739] = 1'd0;
    assign memfont[1740] = 1'd0;
    assign memfont[1741] = 1'd0;
    assign memfont[1742] = 1'd0;
    assign memfont[1743] = 1'd0;
    assign memfont[1744] = 1'd1;
    assign memfont[1745] = 1'd1;
    assign memfont[1746] = 1'd1;
    assign memfont[1747] = 1'd1;
    assign memfont[1748] = 1'd0;
    assign memfont[1749] = 1'd0;
    assign memfont[1750] = 1'd0;
    assign memfont[1751] = 1'd0;
    assign memfont[1752] = 1'd0;
    assign memfont[1753] = 1'd1;
    assign memfont[1754] = 1'd1;
    assign memfont[1755] = 1'd0;
    assign memfont[1756] = 1'd0;
    assign memfont[1757] = 1'd0;
    assign memfont[1758] = 1'd0;
    assign memfont[1759] = 1'd0;
    assign memfont[1760] = 1'd1;
    assign memfont[1761] = 1'd1;
    assign memfont[1762] = 1'd1;
    assign memfont[1763] = 1'd0;
    assign memfont[1764] = 1'd0;
    assign memfont[1765] = 1'd1;
    assign memfont[1766] = 1'd1;
    assign memfont[1767] = 1'd1;
    assign memfont[1768] = 1'd0;
    assign memfont[1769] = 1'd0;
    assign memfont[1770] = 1'd0;
    assign memfont[1771] = 1'd0;
    assign memfont[1772] = 1'd0;
    assign memfont[1773] = 1'd1;
    assign memfont[1774] = 1'd1;
    assign memfont[1775] = 1'd0;
    assign memfont[1776] = 1'd0;
    assign memfont[1777] = 1'd1;
    assign memfont[1778] = 1'd1;
    assign memfont[1779] = 1'd0;
    assign memfont[1780] = 1'd0;
    assign memfont[1781] = 1'd0;
    assign memfont[1782] = 1'd0;
    assign memfont[1783] = 1'd0;
    assign memfont[1784] = 1'd1;
    assign memfont[1785] = 1'd1;
    assign memfont[1786] = 1'd0;
    assign memfont[1787] = 1'd0;
    assign memfont[1788] = 1'd0;
    assign memfont[1789] = 1'd1;
    assign memfont[1790] = 1'd1;
    assign memfont[1791] = 1'd0;
    assign memfont[1792] = 1'd0;
    assign memfont[1793] = 1'd0;
    assign memfont[1794] = 1'd0;
    assign memfont[1795] = 1'd0;
    assign memfont[1796] = 1'd0;
    assign memfont[1797] = 1'd0;
    assign memfont[1798] = 1'd0;
    assign memfont[1799] = 1'd0;
    assign memfont[1800] = 1'd0;
    assign memfont[1801] = 1'd1;
    assign memfont[1802] = 1'd1;
    assign memfont[1803] = 1'd0;
    assign memfont[1804] = 1'd0;
    assign memfont[1805] = 1'd0;
    assign memfont[1806] = 1'd0;
    assign memfont[1807] = 1'd0;
    assign memfont[1808] = 1'd0;
    assign memfont[1809] = 1'd0;
    assign memfont[1810] = 1'd0;
    assign memfont[1811] = 1'd0;
    assign memfont[1812] = 1'd0;
    assign memfont[1813] = 1'd1;
    assign memfont[1814] = 1'd1;
    assign memfont[1815] = 1'd1;
    assign memfont[1816] = 1'd0;
    assign memfont[1817] = 1'd0;
    assign memfont[1818] = 1'd0;
    assign memfont[1819] = 1'd0;
    assign memfont[1820] = 1'd1;
    assign memfont[1821] = 1'd1;
    assign memfont[1822] = 1'd1;
    assign memfont[1823] = 1'd0;
    assign memfont[1824] = 1'd0;
    assign memfont[1825] = 1'd1;
    assign memfont[1826] = 1'd1;
    assign memfont[1827] = 1'd0;
    assign memfont[1828] = 1'd0;
    assign memfont[1829] = 1'd0;
    assign memfont[1830] = 1'd0;
    assign memfont[1831] = 1'd0;
    assign memfont[1832] = 1'd0;
    assign memfont[1833] = 1'd1;
    assign memfont[1834] = 1'd1;
    assign memfont[1835] = 1'd0;
    assign memfont[1836] = 1'd0;
    assign memfont[1837] = 1'd0;
    assign memfont[1838] = 1'd0;
    assign memfont[1839] = 1'd0;
    assign memfont[1840] = 1'd0;
    assign memfont[1841] = 1'd1;
    assign memfont[1842] = 1'd1;
    assign memfont[1843] = 1'd0;
    assign memfont[1844] = 1'd0;
    assign memfont[1845] = 1'd0;
    assign memfont[1846] = 1'd0;
    assign memfont[1847] = 1'd0;
    assign memfont[1848] = 1'd0;
    assign memfont[1849] = 1'd0;
    assign memfont[1850] = 1'd0;
    assign memfont[1851] = 1'd0;
    assign memfont[1852] = 1'd0;
    assign memfont[1853] = 1'd0;
    assign memfont[1854] = 1'd0;
    assign memfont[1855] = 1'd0;
    assign memfont[1856] = 1'd1;
    assign memfont[1857] = 1'd1;
    assign memfont[1858] = 1'd1;
    assign memfont[1859] = 1'd0;
    assign memfont[1860] = 1'd0;
    assign memfont[1861] = 1'd1;
    assign memfont[1862] = 1'd1;
    assign memfont[1863] = 1'd0;
    assign memfont[1864] = 1'd0;
    assign memfont[1865] = 1'd1;
    assign memfont[1866] = 1'd1;
    assign memfont[1867] = 1'd1;
    assign memfont[1868] = 1'd0;
    assign memfont[1869] = 1'd0;
    assign memfont[1870] = 1'd0;
    assign memfont[1871] = 1'd0;
    assign memfont[1872] = 1'd0;
    assign memfont[1873] = 1'd1;
    assign memfont[1874] = 1'd1;
    assign memfont[1875] = 1'd0;
    assign memfont[1876] = 1'd0;
    assign memfont[1877] = 1'd0;
    assign memfont[1878] = 1'd0;
    assign memfont[1879] = 1'd0;
    assign memfont[1880] = 1'd0;
    assign memfont[1881] = 1'd0;
    assign memfont[1882] = 1'd0;
    assign memfont[1883] = 1'd0;
    assign memfont[1884] = 1'd0;
    assign memfont[1885] = 1'd1;
    assign memfont[1886] = 1'd1;
    assign memfont[1887] = 1'd1;
    assign memfont[1888] = 1'd1;
    assign memfont[1889] = 1'd0;
    assign memfont[1890] = 1'd0;
    assign memfont[1891] = 1'd1;
    assign memfont[1892] = 1'd1;
    assign memfont[1893] = 1'd1;
    assign memfont[1894] = 1'd1;
    assign memfont[1895] = 1'd0;
    assign memfont[1896] = 1'd0;
    assign memfont[1897] = 1'd1;
    assign memfont[1898] = 1'd1;
    assign memfont[1899] = 1'd1;
    assign memfont[1900] = 1'd1;
    assign memfont[1901] = 1'd0;
    assign memfont[1902] = 1'd0;
    assign memfont[1903] = 1'd0;
    assign memfont[1904] = 1'd0;
    assign memfont[1905] = 1'd1;
    assign memfont[1906] = 1'd1;
    assign memfont[1907] = 1'd0;
    assign memfont[1908] = 1'd0;
    assign memfont[1909] = 1'd1;
    assign memfont[1910] = 1'd1;
    assign memfont[1911] = 1'd0;
    assign memfont[1912] = 1'd0;
    assign memfont[1913] = 1'd0;
    assign memfont[1914] = 1'd0;
    assign memfont[1915] = 1'd0;
    assign memfont[1916] = 1'd1;
    assign memfont[1917] = 1'd1;
    assign memfont[1918] = 1'd1;
    assign memfont[1919] = 1'd0;
    assign memfont[1920] = 1'd0;
    assign memfont[1921] = 1'd1;
    assign memfont[1922] = 1'd1;
    assign memfont[1923] = 1'd0;
    assign memfont[1924] = 1'd0;
    assign memfont[1925] = 1'd0;
    assign memfont[1926] = 1'd0;
    assign memfont[1927] = 1'd0;
    assign memfont[1928] = 1'd0;
    assign memfont[1929] = 1'd1;
    assign memfont[1930] = 1'd1;
    assign memfont[1931] = 1'd0;
    assign memfont[1932] = 1'd0;
    assign memfont[1933] = 1'd1;
    assign memfont[1934] = 1'd1;
    assign memfont[1935] = 1'd0;
    assign memfont[1936] = 1'd0;
    assign memfont[1937] = 1'd0;
    assign memfont[1938] = 1'd0;
    assign memfont[1939] = 1'd0;
    assign memfont[1940] = 1'd1;
    assign memfont[1941] = 1'd1;
    assign memfont[1942] = 1'd1;
    assign memfont[1943] = 1'd0;
    assign memfont[1944] = 1'd0;
    assign memfont[1945] = 1'd1;
    assign memfont[1946] = 1'd1;
    assign memfont[1947] = 1'd0;
    assign memfont[1948] = 1'd0;
    assign memfont[1949] = 1'd0;
    assign memfont[1950] = 1'd0;
    assign memfont[1951] = 1'd0;
    assign memfont[1952] = 1'd0;
    assign memfont[1953] = 1'd1;
    assign memfont[1954] = 1'd1;
    assign memfont[1955] = 1'd0;
    assign memfont[1956] = 1'd0;
    assign memfont[1957] = 1'd1;
    assign memfont[1958] = 1'd1;
    assign memfont[1959] = 1'd0;
    assign memfont[1960] = 1'd0;
    assign memfont[1961] = 1'd0;
    assign memfont[1962] = 1'd0;
    assign memfont[1963] = 1'd0;
    assign memfont[1964] = 1'd1;
    assign memfont[1965] = 1'd1;
    assign memfont[1966] = 1'd0;
    assign memfont[1967] = 1'd0;
    assign memfont[1968] = 1'd0;
    assign memfont[1969] = 1'd0;
    assign memfont[1970] = 1'd0;
    assign memfont[1971] = 1'd0;
    assign memfont[1972] = 1'd0;
    assign memfont[1973] = 1'd1;
    assign memfont[1974] = 1'd1;
    assign memfont[1975] = 1'd0;
    assign memfont[1976] = 1'd0;
    assign memfont[1977] = 1'd0;
    assign memfont[1978] = 1'd0;
    assign memfont[1979] = 1'd0;
    assign memfont[1980] = 1'd0;
    assign memfont[1981] = 1'd1;
    assign memfont[1982] = 1'd1;
    assign memfont[1983] = 1'd0;
    assign memfont[1984] = 1'd0;
    assign memfont[1985] = 1'd0;
    assign memfont[1986] = 1'd0;
    assign memfont[1987] = 1'd0;
    assign memfont[1988] = 1'd0;
    assign memfont[1989] = 1'd1;
    assign memfont[1990] = 1'd1;
    assign memfont[1991] = 1'd0;
    assign memfont[1992] = 1'd0;
    assign memfont[1993] = 1'd1;
    assign memfont[1994] = 1'd1;
    assign memfont[1995] = 1'd1;
    assign memfont[1996] = 1'd0;
    assign memfont[1997] = 1'd0;
    assign memfont[1998] = 1'd0;
    assign memfont[1999] = 1'd0;
    assign memfont[2000] = 1'd1;
    assign memfont[2001] = 1'd1;
    assign memfont[2002] = 1'd0;
    assign memfont[2003] = 1'd0;
    assign memfont[2004] = 1'd0;
    assign memfont[2005] = 1'd1;
    assign memfont[2006] = 1'd1;
    assign memfont[2007] = 1'd0;
    assign memfont[2008] = 1'd1;
    assign memfont[2009] = 1'd1;
    assign memfont[2010] = 1'd1;
    assign memfont[2011] = 1'd0;
    assign memfont[2012] = 1'd0;
    assign memfont[2013] = 1'd1;
    assign memfont[2014] = 1'd1;
    assign memfont[2015] = 1'd0;
    assign memfont[2016] = 1'd0;
    assign memfont[2017] = 1'd0;
    assign memfont[2018] = 1'd0;
    assign memfont[2019] = 1'd1;
    assign memfont[2020] = 1'd1;
    assign memfont[2021] = 1'd0;
    assign memfont[2022] = 1'd0;
    assign memfont[2023] = 1'd1;
    assign memfont[2024] = 1'd1;
    assign memfont[2025] = 1'd0;
    assign memfont[2026] = 1'd0;
    assign memfont[2027] = 1'd0;
    assign memfont[2028] = 1'd0;
    assign memfont[2029] = 1'd0;
    assign memfont[2030] = 1'd1;
    assign memfont[2031] = 1'd1;
    assign memfont[2032] = 1'd0;
    assign memfont[2033] = 1'd0;
    assign memfont[2034] = 1'd0;
    assign memfont[2035] = 1'd1;
    assign memfont[2036] = 1'd1;
    assign memfont[2037] = 1'd0;
    assign memfont[2038] = 1'd0;
    assign memfont[2039] = 1'd0;
    assign memfont[2040] = 1'd0;
    assign memfont[2041] = 1'd0;
    assign memfont[2042] = 1'd0;
    assign memfont[2043] = 1'd0;
    assign memfont[2044] = 1'd0;
    assign memfont[2045] = 1'd0;
    assign memfont[2046] = 1'd0;
    assign memfont[2047] = 1'd1;
    assign memfont[2048] = 1'd1;
    assign memfont[2049] = 1'd0;
    assign memfont[2050] = 1'd0;
    assign memfont[2051] = 1'd0;
    assign memfont[2052] = 1'd0;
    assign memfont[2053] = 1'd0;
    assign memfont[2054] = 1'd0;
    assign memfont[2055] = 1'd0;
    assign memfont[2056] = 1'd0;
    assign memfont[2057] = 1'd1;
    assign memfont[2058] = 1'd1;
    assign memfont[2059] = 1'd0;
    assign memfont[2060] = 1'd0;
    assign memfont[2061] = 1'd0;
    assign memfont[2062] = 1'd0;
    assign memfont[2063] = 1'd0;
    assign memfont[2064] = 1'd0;
    assign memfont[2065] = 1'd1;
    assign memfont[2066] = 1'd1;
    assign memfont[2067] = 1'd1;
    assign memfont[2068] = 1'd0;
    assign memfont[2069] = 1'd0;
    assign memfont[2070] = 1'd0;
    assign memfont[2071] = 1'd0;
    assign memfont[2072] = 1'd0;
    assign memfont[2073] = 1'd1;
    assign memfont[2074] = 1'd1;
    assign memfont[2075] = 1'd0;
    assign memfont[2076] = 1'd0;
    assign memfont[2077] = 1'd1;
    assign memfont[2078] = 1'd1;
    assign memfont[2079] = 1'd1;
    assign memfont[2080] = 1'd1;
    assign memfont[2081] = 1'd1;
    assign memfont[2082] = 1'd1;
    assign memfont[2083] = 1'd1;
    assign memfont[2084] = 1'd1;
    assign memfont[2085] = 1'd1;
    assign memfont[2086] = 1'd1;
    assign memfont[2087] = 1'd0;
    assign memfont[2088] = 1'd0;
    assign memfont[2089] = 1'd0;
    assign memfont[2090] = 1'd0;
    assign memfont[2091] = 1'd1;
    assign memfont[2092] = 1'd1;
    assign memfont[2093] = 1'd0;
    assign memfont[2094] = 1'd1;
    assign memfont[2095] = 1'd1;
    assign memfont[2096] = 1'd0;
    assign memfont[2097] = 1'd0;
    assign memfont[2098] = 1'd0;
    assign memfont[2099] = 1'd0;
    assign memfont[2100] = 1'd0;
    assign memfont[2101] = 1'd1;
    assign memfont[2102] = 1'd1;
    assign memfont[2103] = 1'd0;
    assign memfont[2104] = 1'd0;
    assign memfont[2105] = 1'd0;
    assign memfont[2106] = 1'd0;
    assign memfont[2107] = 1'd0;
    assign memfont[2108] = 1'd1;
    assign memfont[2109] = 1'd1;
    assign memfont[2110] = 1'd1;
    assign memfont[2111] = 1'd0;
    assign memfont[2112] = 1'd0;
    assign memfont[2113] = 1'd1;
    assign memfont[2114] = 1'd1;
    assign memfont[2115] = 1'd0;
    assign memfont[2116] = 1'd0;
    assign memfont[2117] = 1'd0;
    assign memfont[2118] = 1'd0;
    assign memfont[2119] = 1'd0;
    assign memfont[2120] = 1'd0;
    assign memfont[2121] = 1'd1;
    assign memfont[2122] = 1'd1;
    assign memfont[2123] = 1'd0;
    assign memfont[2124] = 1'd0;
    assign memfont[2125] = 1'd1;
    assign memfont[2126] = 1'd1;
    assign memfont[2127] = 1'd0;
    assign memfont[2128] = 1'd0;
    assign memfont[2129] = 1'd0;
    assign memfont[2130] = 1'd0;
    assign memfont[2131] = 1'd0;
    assign memfont[2132] = 1'd1;
    assign memfont[2133] = 1'd1;
    assign memfont[2134] = 1'd1;
    assign memfont[2135] = 1'd0;
    assign memfont[2136] = 1'd0;
    assign memfont[2137] = 1'd1;
    assign memfont[2138] = 1'd1;
    assign memfont[2139] = 1'd0;
    assign memfont[2140] = 1'd0;
    assign memfont[2141] = 1'd0;
    assign memfont[2142] = 1'd0;
    assign memfont[2143] = 1'd0;
    assign memfont[2144] = 1'd0;
    assign memfont[2145] = 1'd0;
    assign memfont[2146] = 1'd0;
    assign memfont[2147] = 1'd0;
    assign memfont[2148] = 1'd0;
    assign memfont[2149] = 1'd1;
    assign memfont[2150] = 1'd1;
    assign memfont[2151] = 1'd0;
    assign memfont[2152] = 1'd0;
    assign memfont[2153] = 1'd0;
    assign memfont[2154] = 1'd0;
    assign memfont[2155] = 1'd0;
    assign memfont[2156] = 1'd0;
    assign memfont[2157] = 1'd0;
    assign memfont[2158] = 1'd0;
    assign memfont[2159] = 1'd0;
    assign memfont[2160] = 1'd0;
    assign memfont[2161] = 1'd1;
    assign memfont[2162] = 1'd1;
    assign memfont[2163] = 1'd0;
    assign memfont[2164] = 1'd0;
    assign memfont[2165] = 1'd0;
    assign memfont[2166] = 1'd0;
    assign memfont[2167] = 1'd0;
    assign memfont[2168] = 1'd0;
    assign memfont[2169] = 1'd1;
    assign memfont[2170] = 1'd1;
    assign memfont[2171] = 1'd0;
    assign memfont[2172] = 1'd0;
    assign memfont[2173] = 1'd1;
    assign memfont[2174] = 1'd1;
    assign memfont[2175] = 1'd0;
    assign memfont[2176] = 1'd0;
    assign memfont[2177] = 1'd0;
    assign memfont[2178] = 1'd0;
    assign memfont[2179] = 1'd0;
    assign memfont[2180] = 1'd0;
    assign memfont[2181] = 1'd1;
    assign memfont[2182] = 1'd1;
    assign memfont[2183] = 1'd0;
    assign memfont[2184] = 1'd0;
    assign memfont[2185] = 1'd0;
    assign memfont[2186] = 1'd0;
    assign memfont[2187] = 1'd0;
    assign memfont[2188] = 1'd0;
    assign memfont[2189] = 1'd1;
    assign memfont[2190] = 1'd1;
    assign memfont[2191] = 1'd0;
    assign memfont[2192] = 1'd0;
    assign memfont[2193] = 1'd0;
    assign memfont[2194] = 1'd0;
    assign memfont[2195] = 1'd0;
    assign memfont[2196] = 1'd0;
    assign memfont[2197] = 1'd0;
    assign memfont[2198] = 1'd0;
    assign memfont[2199] = 1'd0;
    assign memfont[2200] = 1'd0;
    assign memfont[2201] = 1'd0;
    assign memfont[2202] = 1'd0;
    assign memfont[2203] = 1'd0;
    assign memfont[2204] = 1'd1;
    assign memfont[2205] = 1'd1;
    assign memfont[2206] = 1'd1;
    assign memfont[2207] = 1'd0;
    assign memfont[2208] = 1'd0;
    assign memfont[2209] = 1'd1;
    assign memfont[2210] = 1'd1;
    assign memfont[2211] = 1'd0;
    assign memfont[2212] = 1'd0;
    assign memfont[2213] = 1'd1;
    assign memfont[2214] = 1'd1;
    assign memfont[2215] = 1'd0;
    assign memfont[2216] = 1'd0;
    assign memfont[2217] = 1'd0;
    assign memfont[2218] = 1'd0;
    assign memfont[2219] = 1'd0;
    assign memfont[2220] = 1'd0;
    assign memfont[2221] = 1'd1;
    assign memfont[2222] = 1'd1;
    assign memfont[2223] = 1'd0;
    assign memfont[2224] = 1'd0;
    assign memfont[2225] = 1'd0;
    assign memfont[2226] = 1'd0;
    assign memfont[2227] = 1'd0;
    assign memfont[2228] = 1'd0;
    assign memfont[2229] = 1'd0;
    assign memfont[2230] = 1'd0;
    assign memfont[2231] = 1'd0;
    assign memfont[2232] = 1'd0;
    assign memfont[2233] = 1'd1;
    assign memfont[2234] = 1'd1;
    assign memfont[2235] = 1'd1;
    assign memfont[2236] = 1'd1;
    assign memfont[2237] = 1'd0;
    assign memfont[2238] = 1'd0;
    assign memfont[2239] = 1'd1;
    assign memfont[2240] = 1'd1;
    assign memfont[2241] = 1'd1;
    assign memfont[2242] = 1'd1;
    assign memfont[2243] = 1'd0;
    assign memfont[2244] = 1'd0;
    assign memfont[2245] = 1'd1;
    assign memfont[2246] = 1'd1;
    assign memfont[2247] = 1'd1;
    assign memfont[2248] = 1'd1;
    assign memfont[2249] = 1'd0;
    assign memfont[2250] = 1'd0;
    assign memfont[2251] = 1'd0;
    assign memfont[2252] = 1'd0;
    assign memfont[2253] = 1'd1;
    assign memfont[2254] = 1'd1;
    assign memfont[2255] = 1'd0;
    assign memfont[2256] = 1'd0;
    assign memfont[2257] = 1'd1;
    assign memfont[2258] = 1'd1;
    assign memfont[2259] = 1'd0;
    assign memfont[2260] = 1'd0;
    assign memfont[2261] = 1'd0;
    assign memfont[2262] = 1'd0;
    assign memfont[2263] = 1'd0;
    assign memfont[2264] = 1'd0;
    assign memfont[2265] = 1'd1;
    assign memfont[2266] = 1'd1;
    assign memfont[2267] = 1'd0;
    assign memfont[2268] = 1'd0;
    assign memfont[2269] = 1'd1;
    assign memfont[2270] = 1'd1;
    assign memfont[2271] = 1'd0;
    assign memfont[2272] = 1'd0;
    assign memfont[2273] = 1'd0;
    assign memfont[2274] = 1'd0;
    assign memfont[2275] = 1'd0;
    assign memfont[2276] = 1'd0;
    assign memfont[2277] = 1'd1;
    assign memfont[2278] = 1'd1;
    assign memfont[2279] = 1'd0;
    assign memfont[2280] = 1'd0;
    assign memfont[2281] = 1'd1;
    assign memfont[2282] = 1'd1;
    assign memfont[2283] = 1'd0;
    assign memfont[2284] = 1'd0;
    assign memfont[2285] = 1'd0;
    assign memfont[2286] = 1'd0;
    assign memfont[2287] = 1'd0;
    assign memfont[2288] = 1'd0;
    assign memfont[2289] = 1'd1;
    assign memfont[2290] = 1'd1;
    assign memfont[2291] = 1'd0;
    assign memfont[2292] = 1'd0;
    assign memfont[2293] = 1'd1;
    assign memfont[2294] = 1'd1;
    assign memfont[2295] = 1'd0;
    assign memfont[2296] = 1'd0;
    assign memfont[2297] = 1'd0;
    assign memfont[2298] = 1'd0;
    assign memfont[2299] = 1'd0;
    assign memfont[2300] = 1'd0;
    assign memfont[2301] = 1'd1;
    assign memfont[2302] = 1'd1;
    assign memfont[2303] = 1'd0;
    assign memfont[2304] = 1'd0;
    assign memfont[2305] = 1'd1;
    assign memfont[2306] = 1'd1;
    assign memfont[2307] = 1'd1;
    assign memfont[2308] = 1'd0;
    assign memfont[2309] = 1'd0;
    assign memfont[2310] = 1'd0;
    assign memfont[2311] = 1'd0;
    assign memfont[2312] = 1'd0;
    assign memfont[2313] = 1'd0;
    assign memfont[2314] = 1'd0;
    assign memfont[2315] = 1'd0;
    assign memfont[2316] = 1'd0;
    assign memfont[2317] = 1'd0;
    assign memfont[2318] = 1'd0;
    assign memfont[2319] = 1'd0;
    assign memfont[2320] = 1'd0;
    assign memfont[2321] = 1'd1;
    assign memfont[2322] = 1'd1;
    assign memfont[2323] = 1'd0;
    assign memfont[2324] = 1'd0;
    assign memfont[2325] = 1'd0;
    assign memfont[2326] = 1'd0;
    assign memfont[2327] = 1'd0;
    assign memfont[2328] = 1'd0;
    assign memfont[2329] = 1'd1;
    assign memfont[2330] = 1'd1;
    assign memfont[2331] = 1'd0;
    assign memfont[2332] = 1'd0;
    assign memfont[2333] = 1'd0;
    assign memfont[2334] = 1'd0;
    assign memfont[2335] = 1'd0;
    assign memfont[2336] = 1'd0;
    assign memfont[2337] = 1'd1;
    assign memfont[2338] = 1'd1;
    assign memfont[2339] = 1'd0;
    assign memfont[2340] = 1'd0;
    assign memfont[2341] = 1'd0;
    assign memfont[2342] = 1'd1;
    assign memfont[2343] = 1'd1;
    assign memfont[2344] = 1'd0;
    assign memfont[2345] = 1'd0;
    assign memfont[2346] = 1'd0;
    assign memfont[2347] = 1'd0;
    assign memfont[2348] = 1'd1;
    assign memfont[2349] = 1'd1;
    assign memfont[2350] = 1'd0;
    assign memfont[2351] = 1'd0;
    assign memfont[2352] = 1'd0;
    assign memfont[2353] = 1'd1;
    assign memfont[2354] = 1'd1;
    assign memfont[2355] = 1'd0;
    assign memfont[2356] = 1'd1;
    assign memfont[2357] = 1'd1;
    assign memfont[2358] = 1'd1;
    assign memfont[2359] = 1'd1;
    assign memfont[2360] = 1'd0;
    assign memfont[2361] = 1'd1;
    assign memfont[2362] = 1'd1;
    assign memfont[2363] = 1'd0;
    assign memfont[2364] = 1'd0;
    assign memfont[2365] = 1'd0;
    assign memfont[2366] = 1'd0;
    assign memfont[2367] = 1'd1;
    assign memfont[2368] = 1'd1;
    assign memfont[2369] = 1'd0;
    assign memfont[2370] = 1'd1;
    assign memfont[2371] = 1'd1;
    assign memfont[2372] = 1'd0;
    assign memfont[2373] = 1'd0;
    assign memfont[2374] = 1'd0;
    assign memfont[2375] = 1'd0;
    assign memfont[2376] = 1'd0;
    assign memfont[2377] = 1'd0;
    assign memfont[2378] = 1'd0;
    assign memfont[2379] = 1'd1;
    assign memfont[2380] = 1'd1;
    assign memfont[2381] = 1'd0;
    assign memfont[2382] = 1'd0;
    assign memfont[2383] = 1'd1;
    assign memfont[2384] = 1'd1;
    assign memfont[2385] = 1'd0;
    assign memfont[2386] = 1'd0;
    assign memfont[2387] = 1'd0;
    assign memfont[2388] = 1'd0;
    assign memfont[2389] = 1'd0;
    assign memfont[2390] = 1'd0;
    assign memfont[2391] = 1'd0;
    assign memfont[2392] = 1'd0;
    assign memfont[2393] = 1'd0;
    assign memfont[2394] = 1'd1;
    assign memfont[2395] = 1'd1;
    assign memfont[2396] = 1'd1;
    assign memfont[2397] = 1'd0;
    assign memfont[2398] = 1'd0;
    assign memfont[2399] = 1'd0;
    assign memfont[2400] = 1'd0;
    assign memfont[2401] = 1'd0;
    assign memfont[2402] = 1'd0;
    assign memfont[2403] = 1'd0;
    assign memfont[2404] = 1'd0;
    assign memfont[2405] = 1'd1;
    assign memfont[2406] = 1'd1;
    assign memfont[2407] = 1'd0;
    assign memfont[2408] = 1'd0;
    assign memfont[2409] = 1'd0;
    assign memfont[2410] = 1'd0;
    assign memfont[2411] = 1'd0;
    assign memfont[2412] = 1'd0;
    assign memfont[2413] = 1'd1;
    assign memfont[2414] = 1'd1;
    assign memfont[2415] = 1'd1;
    assign memfont[2416] = 1'd0;
    assign memfont[2417] = 1'd0;
    assign memfont[2418] = 1'd1;
    assign memfont[2419] = 1'd1;
    assign memfont[2420] = 1'd1;
    assign memfont[2421] = 1'd1;
    assign memfont[2422] = 1'd1;
    assign memfont[2423] = 1'd0;
    assign memfont[2424] = 1'd0;
    assign memfont[2425] = 1'd1;
    assign memfont[2426] = 1'd1;
    assign memfont[2427] = 1'd1;
    assign memfont[2428] = 1'd1;
    assign memfont[2429] = 1'd0;
    assign memfont[2430] = 1'd0;
    assign memfont[2431] = 1'd1;
    assign memfont[2432] = 1'd1;
    assign memfont[2433] = 1'd1;
    assign memfont[2434] = 1'd1;
    assign memfont[2435] = 1'd0;
    assign memfont[2436] = 1'd0;
    assign memfont[2437] = 1'd0;
    assign memfont[2438] = 1'd0;
    assign memfont[2439] = 1'd1;
    assign memfont[2440] = 1'd1;
    assign memfont[2441] = 1'd0;
    assign memfont[2442] = 1'd0;
    assign memfont[2443] = 1'd1;
    assign memfont[2444] = 1'd1;
    assign memfont[2445] = 1'd0;
    assign memfont[2446] = 1'd0;
    assign memfont[2447] = 1'd0;
    assign memfont[2448] = 1'd0;
    assign memfont[2449] = 1'd1;
    assign memfont[2450] = 1'd1;
    assign memfont[2451] = 1'd0;
    assign memfont[2452] = 1'd0;
    assign memfont[2453] = 1'd0;
    assign memfont[2454] = 1'd0;
    assign memfont[2455] = 1'd0;
    assign memfont[2456] = 1'd1;
    assign memfont[2457] = 1'd1;
    assign memfont[2458] = 1'd0;
    assign memfont[2459] = 1'd0;
    assign memfont[2460] = 1'd0;
    assign memfont[2461] = 1'd1;
    assign memfont[2462] = 1'd1;
    assign memfont[2463] = 1'd0;
    assign memfont[2464] = 1'd0;
    assign memfont[2465] = 1'd0;
    assign memfont[2466] = 1'd0;
    assign memfont[2467] = 1'd0;
    assign memfont[2468] = 1'd0;
    assign memfont[2469] = 1'd0;
    assign memfont[2470] = 1'd0;
    assign memfont[2471] = 1'd0;
    assign memfont[2472] = 1'd0;
    assign memfont[2473] = 1'd1;
    assign memfont[2474] = 1'd1;
    assign memfont[2475] = 1'd0;
    assign memfont[2476] = 1'd0;
    assign memfont[2477] = 1'd0;
    assign memfont[2478] = 1'd0;
    assign memfont[2479] = 1'd0;
    assign memfont[2480] = 1'd0;
    assign memfont[2481] = 1'd1;
    assign memfont[2482] = 1'd1;
    assign memfont[2483] = 1'd0;
    assign memfont[2484] = 1'd0;
    assign memfont[2485] = 1'd1;
    assign memfont[2486] = 1'd1;
    assign memfont[2487] = 1'd0;
    assign memfont[2488] = 1'd0;
    assign memfont[2489] = 1'd0;
    assign memfont[2490] = 1'd0;
    assign memfont[2491] = 1'd0;
    assign memfont[2492] = 1'd0;
    assign memfont[2493] = 1'd0;
    assign memfont[2494] = 1'd0;
    assign memfont[2495] = 1'd0;
    assign memfont[2496] = 1'd0;
    assign memfont[2497] = 1'd1;
    assign memfont[2498] = 1'd1;
    assign memfont[2499] = 1'd0;
    assign memfont[2500] = 1'd0;
    assign memfont[2501] = 1'd0;
    assign memfont[2502] = 1'd0;
    assign memfont[2503] = 1'd0;
    assign memfont[2504] = 1'd0;
    assign memfont[2505] = 1'd0;
    assign memfont[2506] = 1'd0;
    assign memfont[2507] = 1'd0;
    assign memfont[2508] = 1'd0;
    assign memfont[2509] = 1'd1;
    assign memfont[2510] = 1'd1;
    assign memfont[2511] = 1'd0;
    assign memfont[2512] = 1'd0;
    assign memfont[2513] = 1'd0;
    assign memfont[2514] = 1'd0;
    assign memfont[2515] = 1'd0;
    assign memfont[2516] = 1'd0;
    assign memfont[2517] = 1'd0;
    assign memfont[2518] = 1'd0;
    assign memfont[2519] = 1'd0;
    assign memfont[2520] = 1'd0;
    assign memfont[2521] = 1'd1;
    assign memfont[2522] = 1'd1;
    assign memfont[2523] = 1'd0;
    assign memfont[2524] = 1'd0;
    assign memfont[2525] = 1'd0;
    assign memfont[2526] = 1'd0;
    assign memfont[2527] = 1'd0;
    assign memfont[2528] = 1'd0;
    assign memfont[2529] = 1'd1;
    assign memfont[2530] = 1'd1;
    assign memfont[2531] = 1'd0;
    assign memfont[2532] = 1'd0;
    assign memfont[2533] = 1'd0;
    assign memfont[2534] = 1'd0;
    assign memfont[2535] = 1'd0;
    assign memfont[2536] = 1'd0;
    assign memfont[2537] = 1'd1;
    assign memfont[2538] = 1'd1;
    assign memfont[2539] = 1'd0;
    assign memfont[2540] = 1'd0;
    assign memfont[2541] = 1'd0;
    assign memfont[2542] = 1'd0;
    assign memfont[2543] = 1'd0;
    assign memfont[2544] = 1'd0;
    assign memfont[2545] = 1'd0;
    assign memfont[2546] = 1'd0;
    assign memfont[2547] = 1'd0;
    assign memfont[2548] = 1'd0;
    assign memfont[2549] = 1'd0;
    assign memfont[2550] = 1'd0;
    assign memfont[2551] = 1'd0;
    assign memfont[2552] = 1'd1;
    assign memfont[2553] = 1'd1;
    assign memfont[2554] = 1'd1;
    assign memfont[2555] = 1'd0;
    assign memfont[2556] = 1'd0;
    assign memfont[2557] = 1'd1;
    assign memfont[2558] = 1'd1;
    assign memfont[2559] = 1'd0;
    assign memfont[2560] = 1'd1;
    assign memfont[2561] = 1'd1;
    assign memfont[2562] = 1'd0;
    assign memfont[2563] = 1'd0;
    assign memfont[2564] = 1'd0;
    assign memfont[2565] = 1'd0;
    assign memfont[2566] = 1'd0;
    assign memfont[2567] = 1'd0;
    assign memfont[2568] = 1'd0;
    assign memfont[2569] = 1'd1;
    assign memfont[2570] = 1'd1;
    assign memfont[2571] = 1'd0;
    assign memfont[2572] = 1'd0;
    assign memfont[2573] = 1'd0;
    assign memfont[2574] = 1'd0;
    assign memfont[2575] = 1'd0;
    assign memfont[2576] = 1'd0;
    assign memfont[2577] = 1'd0;
    assign memfont[2578] = 1'd0;
    assign memfont[2579] = 1'd0;
    assign memfont[2580] = 1'd0;
    assign memfont[2581] = 1'd1;
    assign memfont[2582] = 1'd1;
    assign memfont[2583] = 1'd1;
    assign memfont[2584] = 1'd1;
    assign memfont[2585] = 1'd0;
    assign memfont[2586] = 1'd0;
    assign memfont[2587] = 1'd1;
    assign memfont[2588] = 1'd1;
    assign memfont[2589] = 1'd1;
    assign memfont[2590] = 1'd1;
    assign memfont[2591] = 1'd0;
    assign memfont[2592] = 1'd0;
    assign memfont[2593] = 1'd1;
    assign memfont[2594] = 1'd1;
    assign memfont[2595] = 1'd0;
    assign memfont[2596] = 1'd1;
    assign memfont[2597] = 1'd1;
    assign memfont[2598] = 1'd0;
    assign memfont[2599] = 1'd0;
    assign memfont[2600] = 1'd0;
    assign memfont[2601] = 1'd1;
    assign memfont[2602] = 1'd1;
    assign memfont[2603] = 1'd0;
    assign memfont[2604] = 1'd0;
    assign memfont[2605] = 1'd1;
    assign memfont[2606] = 1'd1;
    assign memfont[2607] = 1'd0;
    assign memfont[2608] = 1'd0;
    assign memfont[2609] = 1'd0;
    assign memfont[2610] = 1'd0;
    assign memfont[2611] = 1'd0;
    assign memfont[2612] = 1'd0;
    assign memfont[2613] = 1'd1;
    assign memfont[2614] = 1'd1;
    assign memfont[2615] = 1'd0;
    assign memfont[2616] = 1'd0;
    assign memfont[2617] = 1'd1;
    assign memfont[2618] = 1'd1;
    assign memfont[2619] = 1'd0;
    assign memfont[2620] = 1'd0;
    assign memfont[2621] = 1'd0;
    assign memfont[2622] = 1'd0;
    assign memfont[2623] = 1'd0;
    assign memfont[2624] = 1'd0;
    assign memfont[2625] = 1'd1;
    assign memfont[2626] = 1'd1;
    assign memfont[2627] = 1'd0;
    assign memfont[2628] = 1'd0;
    assign memfont[2629] = 1'd1;
    assign memfont[2630] = 1'd1;
    assign memfont[2631] = 1'd0;
    assign memfont[2632] = 1'd0;
    assign memfont[2633] = 1'd0;
    assign memfont[2634] = 1'd0;
    assign memfont[2635] = 1'd0;
    assign memfont[2636] = 1'd0;
    assign memfont[2637] = 1'd1;
    assign memfont[2638] = 1'd1;
    assign memfont[2639] = 1'd0;
    assign memfont[2640] = 1'd0;
    assign memfont[2641] = 1'd1;
    assign memfont[2642] = 1'd1;
    assign memfont[2643] = 1'd0;
    assign memfont[2644] = 1'd0;
    assign memfont[2645] = 1'd0;
    assign memfont[2646] = 1'd0;
    assign memfont[2647] = 1'd0;
    assign memfont[2648] = 1'd1;
    assign memfont[2649] = 1'd1;
    assign memfont[2650] = 1'd1;
    assign memfont[2651] = 1'd0;
    assign memfont[2652] = 1'd0;
    assign memfont[2653] = 1'd0;
    assign memfont[2654] = 1'd1;
    assign memfont[2655] = 1'd1;
    assign memfont[2656] = 1'd1;
    assign memfont[2657] = 1'd0;
    assign memfont[2658] = 1'd0;
    assign memfont[2659] = 1'd0;
    assign memfont[2660] = 1'd0;
    assign memfont[2661] = 1'd0;
    assign memfont[2662] = 1'd0;
    assign memfont[2663] = 1'd0;
    assign memfont[2664] = 1'd0;
    assign memfont[2665] = 1'd0;
    assign memfont[2666] = 1'd0;
    assign memfont[2667] = 1'd0;
    assign memfont[2668] = 1'd0;
    assign memfont[2669] = 1'd1;
    assign memfont[2670] = 1'd1;
    assign memfont[2671] = 1'd0;
    assign memfont[2672] = 1'd0;
    assign memfont[2673] = 1'd0;
    assign memfont[2674] = 1'd0;
    assign memfont[2675] = 1'd0;
    assign memfont[2676] = 1'd0;
    assign memfont[2677] = 1'd1;
    assign memfont[2678] = 1'd1;
    assign memfont[2679] = 1'd0;
    assign memfont[2680] = 1'd0;
    assign memfont[2681] = 1'd0;
    assign memfont[2682] = 1'd0;
    assign memfont[2683] = 1'd0;
    assign memfont[2684] = 1'd0;
    assign memfont[2685] = 1'd1;
    assign memfont[2686] = 1'd1;
    assign memfont[2687] = 1'd0;
    assign memfont[2688] = 1'd0;
    assign memfont[2689] = 1'd0;
    assign memfont[2690] = 1'd1;
    assign memfont[2691] = 1'd1;
    assign memfont[2692] = 1'd0;
    assign memfont[2693] = 1'd0;
    assign memfont[2694] = 1'd0;
    assign memfont[2695] = 1'd0;
    assign memfont[2696] = 1'd1;
    assign memfont[2697] = 1'd1;
    assign memfont[2698] = 1'd0;
    assign memfont[2699] = 1'd0;
    assign memfont[2700] = 1'd0;
    assign memfont[2701] = 1'd1;
    assign memfont[2702] = 1'd1;
    assign memfont[2703] = 1'd0;
    assign memfont[2704] = 1'd1;
    assign memfont[2705] = 1'd0;
    assign memfont[2706] = 1'd1;
    assign memfont[2707] = 1'd1;
    assign memfont[2708] = 1'd0;
    assign memfont[2709] = 1'd1;
    assign memfont[2710] = 1'd1;
    assign memfont[2711] = 1'd0;
    assign memfont[2712] = 1'd0;
    assign memfont[2713] = 1'd0;
    assign memfont[2714] = 1'd0;
    assign memfont[2715] = 1'd0;
    assign memfont[2716] = 1'd1;
    assign memfont[2717] = 1'd1;
    assign memfont[2718] = 1'd1;
    assign memfont[2719] = 1'd1;
    assign memfont[2720] = 1'd0;
    assign memfont[2721] = 1'd0;
    assign memfont[2722] = 1'd0;
    assign memfont[2723] = 1'd0;
    assign memfont[2724] = 1'd0;
    assign memfont[2725] = 1'd0;
    assign memfont[2726] = 1'd0;
    assign memfont[2727] = 1'd1;
    assign memfont[2728] = 1'd1;
    assign memfont[2729] = 1'd0;
    assign memfont[2730] = 1'd1;
    assign memfont[2731] = 1'd1;
    assign memfont[2732] = 1'd0;
    assign memfont[2733] = 1'd0;
    assign memfont[2734] = 1'd0;
    assign memfont[2735] = 1'd0;
    assign memfont[2736] = 1'd0;
    assign memfont[2737] = 1'd0;
    assign memfont[2738] = 1'd0;
    assign memfont[2739] = 1'd0;
    assign memfont[2740] = 1'd0;
    assign memfont[2741] = 1'd0;
    assign memfont[2742] = 1'd1;
    assign memfont[2743] = 1'd1;
    assign memfont[2744] = 1'd0;
    assign memfont[2745] = 1'd0;
    assign memfont[2746] = 1'd0;
    assign memfont[2747] = 1'd0;
    assign memfont[2748] = 1'd0;
    assign memfont[2749] = 1'd0;
    assign memfont[2750] = 1'd0;
    assign memfont[2751] = 1'd0;
    assign memfont[2752] = 1'd0;
    assign memfont[2753] = 1'd1;
    assign memfont[2754] = 1'd1;
    assign memfont[2755] = 1'd0;
    assign memfont[2756] = 1'd0;
    assign memfont[2757] = 1'd0;
    assign memfont[2758] = 1'd0;
    assign memfont[2759] = 1'd0;
    assign memfont[2760] = 1'd0;
    assign memfont[2761] = 1'd1;
    assign memfont[2762] = 1'd1;
    assign memfont[2763] = 1'd0;
    assign memfont[2764] = 1'd0;
    assign memfont[2765] = 1'd0;
    assign memfont[2766] = 1'd0;
    assign memfont[2767] = 1'd0;
    assign memfont[2768] = 1'd1;
    assign memfont[2769] = 1'd1;
    assign memfont[2770] = 1'd1;
    assign memfont[2771] = 1'd0;
    assign memfont[2772] = 1'd0;
    assign memfont[2773] = 1'd1;
    assign memfont[2774] = 1'd1;
    assign memfont[2775] = 1'd1;
    assign memfont[2776] = 1'd1;
    assign memfont[2777] = 1'd0;
    assign memfont[2778] = 1'd0;
    assign memfont[2779] = 1'd1;
    assign memfont[2780] = 1'd1;
    assign memfont[2781] = 1'd1;
    assign memfont[2782] = 1'd1;
    assign memfont[2783] = 1'd0;
    assign memfont[2784] = 1'd0;
    assign memfont[2785] = 1'd0;
    assign memfont[2786] = 1'd0;
    assign memfont[2787] = 1'd1;
    assign memfont[2788] = 1'd1;
    assign memfont[2789] = 1'd0;
    assign memfont[2790] = 1'd0;
    assign memfont[2791] = 1'd1;
    assign memfont[2792] = 1'd1;
    assign memfont[2793] = 1'd0;
    assign memfont[2794] = 1'd0;
    assign memfont[2795] = 1'd0;
    assign memfont[2796] = 1'd0;
    assign memfont[2797] = 1'd1;
    assign memfont[2798] = 1'd1;
    assign memfont[2799] = 1'd1;
    assign memfont[2800] = 1'd1;
    assign memfont[2801] = 1'd1;
    assign memfont[2802] = 1'd1;
    assign memfont[2803] = 1'd1;
    assign memfont[2804] = 1'd1;
    assign memfont[2805] = 1'd0;
    assign memfont[2806] = 1'd0;
    assign memfont[2807] = 1'd0;
    assign memfont[2808] = 1'd0;
    assign memfont[2809] = 1'd1;
    assign memfont[2810] = 1'd1;
    assign memfont[2811] = 1'd0;
    assign memfont[2812] = 1'd0;
    assign memfont[2813] = 1'd0;
    assign memfont[2814] = 1'd0;
    assign memfont[2815] = 1'd0;
    assign memfont[2816] = 1'd0;
    assign memfont[2817] = 1'd0;
    assign memfont[2818] = 1'd0;
    assign memfont[2819] = 1'd0;
    assign memfont[2820] = 1'd0;
    assign memfont[2821] = 1'd1;
    assign memfont[2822] = 1'd1;
    assign memfont[2823] = 1'd0;
    assign memfont[2824] = 1'd0;
    assign memfont[2825] = 1'd0;
    assign memfont[2826] = 1'd0;
    assign memfont[2827] = 1'd0;
    assign memfont[2828] = 1'd0;
    assign memfont[2829] = 1'd1;
    assign memfont[2830] = 1'd1;
    assign memfont[2831] = 1'd0;
    assign memfont[2832] = 1'd0;
    assign memfont[2833] = 1'd1;
    assign memfont[2834] = 1'd1;
    assign memfont[2835] = 1'd1;
    assign memfont[2836] = 1'd1;
    assign memfont[2837] = 1'd1;
    assign memfont[2838] = 1'd1;
    assign memfont[2839] = 1'd1;
    assign memfont[2840] = 1'd1;
    assign memfont[2841] = 1'd1;
    assign memfont[2842] = 1'd0;
    assign memfont[2843] = 1'd0;
    assign memfont[2844] = 1'd0;
    assign memfont[2845] = 1'd1;
    assign memfont[2846] = 1'd1;
    assign memfont[2847] = 1'd0;
    assign memfont[2848] = 1'd0;
    assign memfont[2849] = 1'd0;
    assign memfont[2850] = 1'd0;
    assign memfont[2851] = 1'd0;
    assign memfont[2852] = 1'd0;
    assign memfont[2853] = 1'd0;
    assign memfont[2854] = 1'd0;
    assign memfont[2855] = 1'd0;
    assign memfont[2856] = 1'd0;
    assign memfont[2857] = 1'd1;
    assign memfont[2858] = 1'd1;
    assign memfont[2859] = 1'd0;
    assign memfont[2860] = 1'd0;
    assign memfont[2861] = 1'd0;
    assign memfont[2862] = 1'd0;
    assign memfont[2863] = 1'd0;
    assign memfont[2864] = 1'd0;
    assign memfont[2865] = 1'd0;
    assign memfont[2866] = 1'd0;
    assign memfont[2867] = 1'd0;
    assign memfont[2868] = 1'd0;
    assign memfont[2869] = 1'd1;
    assign memfont[2870] = 1'd1;
    assign memfont[2871] = 1'd1;
    assign memfont[2872] = 1'd1;
    assign memfont[2873] = 1'd1;
    assign memfont[2874] = 1'd1;
    assign memfont[2875] = 1'd1;
    assign memfont[2876] = 1'd1;
    assign memfont[2877] = 1'd1;
    assign memfont[2878] = 1'd1;
    assign memfont[2879] = 1'd0;
    assign memfont[2880] = 1'd0;
    assign memfont[2881] = 1'd0;
    assign memfont[2882] = 1'd0;
    assign memfont[2883] = 1'd0;
    assign memfont[2884] = 1'd0;
    assign memfont[2885] = 1'd1;
    assign memfont[2886] = 1'd1;
    assign memfont[2887] = 1'd0;
    assign memfont[2888] = 1'd0;
    assign memfont[2889] = 1'd0;
    assign memfont[2890] = 1'd0;
    assign memfont[2891] = 1'd0;
    assign memfont[2892] = 1'd0;
    assign memfont[2893] = 1'd0;
    assign memfont[2894] = 1'd0;
    assign memfont[2895] = 1'd0;
    assign memfont[2896] = 1'd0;
    assign memfont[2897] = 1'd0;
    assign memfont[2898] = 1'd0;
    assign memfont[2899] = 1'd0;
    assign memfont[2900] = 1'd1;
    assign memfont[2901] = 1'd1;
    assign memfont[2902] = 1'd1;
    assign memfont[2903] = 1'd0;
    assign memfont[2904] = 1'd0;
    assign memfont[2905] = 1'd1;
    assign memfont[2906] = 1'd1;
    assign memfont[2907] = 1'd1;
    assign memfont[2908] = 1'd1;
    assign memfont[2909] = 1'd1;
    assign memfont[2910] = 1'd0;
    assign memfont[2911] = 1'd0;
    assign memfont[2912] = 1'd0;
    assign memfont[2913] = 1'd0;
    assign memfont[2914] = 1'd0;
    assign memfont[2915] = 1'd0;
    assign memfont[2916] = 1'd0;
    assign memfont[2917] = 1'd1;
    assign memfont[2918] = 1'd1;
    assign memfont[2919] = 1'd0;
    assign memfont[2920] = 1'd0;
    assign memfont[2921] = 1'd0;
    assign memfont[2922] = 1'd0;
    assign memfont[2923] = 1'd0;
    assign memfont[2924] = 1'd0;
    assign memfont[2925] = 1'd0;
    assign memfont[2926] = 1'd0;
    assign memfont[2927] = 1'd0;
    assign memfont[2928] = 1'd0;
    assign memfont[2929] = 1'd1;
    assign memfont[2930] = 1'd1;
    assign memfont[2931] = 1'd1;
    assign memfont[2932] = 1'd1;
    assign memfont[2933] = 1'd0;
    assign memfont[2934] = 1'd0;
    assign memfont[2935] = 1'd1;
    assign memfont[2936] = 1'd0;
    assign memfont[2937] = 1'd1;
    assign memfont[2938] = 1'd1;
    assign memfont[2939] = 1'd0;
    assign memfont[2940] = 1'd0;
    assign memfont[2941] = 1'd1;
    assign memfont[2942] = 1'd1;
    assign memfont[2943] = 1'd0;
    assign memfont[2944] = 1'd1;
    assign memfont[2945] = 1'd1;
    assign memfont[2946] = 1'd0;
    assign memfont[2947] = 1'd0;
    assign memfont[2948] = 1'd0;
    assign memfont[2949] = 1'd1;
    assign memfont[2950] = 1'd1;
    assign memfont[2951] = 1'd0;
    assign memfont[2952] = 1'd0;
    assign memfont[2953] = 1'd1;
    assign memfont[2954] = 1'd1;
    assign memfont[2955] = 1'd0;
    assign memfont[2956] = 1'd0;
    assign memfont[2957] = 1'd0;
    assign memfont[2958] = 1'd0;
    assign memfont[2959] = 1'd0;
    assign memfont[2960] = 1'd0;
    assign memfont[2961] = 1'd1;
    assign memfont[2962] = 1'd1;
    assign memfont[2963] = 1'd0;
    assign memfont[2964] = 1'd0;
    assign memfont[2965] = 1'd1;
    assign memfont[2966] = 1'd1;
    assign memfont[2967] = 1'd0;
    assign memfont[2968] = 1'd0;
    assign memfont[2969] = 1'd0;
    assign memfont[2970] = 1'd0;
    assign memfont[2971] = 1'd0;
    assign memfont[2972] = 1'd1;
    assign memfont[2973] = 1'd1;
    assign memfont[2974] = 1'd1;
    assign memfont[2975] = 1'd0;
    assign memfont[2976] = 1'd0;
    assign memfont[2977] = 1'd1;
    assign memfont[2978] = 1'd1;
    assign memfont[2979] = 1'd0;
    assign memfont[2980] = 1'd0;
    assign memfont[2981] = 1'd0;
    assign memfont[2982] = 1'd0;
    assign memfont[2983] = 1'd0;
    assign memfont[2984] = 1'd0;
    assign memfont[2985] = 1'd1;
    assign memfont[2986] = 1'd1;
    assign memfont[2987] = 1'd0;
    assign memfont[2988] = 1'd0;
    assign memfont[2989] = 1'd1;
    assign memfont[2990] = 1'd1;
    assign memfont[2991] = 1'd0;
    assign memfont[2992] = 1'd0;
    assign memfont[2993] = 1'd0;
    assign memfont[2994] = 1'd0;
    assign memfont[2995] = 1'd1;
    assign memfont[2996] = 1'd1;
    assign memfont[2997] = 1'd1;
    assign memfont[2998] = 1'd0;
    assign memfont[2999] = 1'd0;
    assign memfont[3000] = 1'd0;
    assign memfont[3001] = 1'd0;
    assign memfont[3002] = 1'd0;
    assign memfont[3003] = 1'd1;
    assign memfont[3004] = 1'd1;
    assign memfont[3005] = 1'd1;
    assign memfont[3006] = 1'd1;
    assign memfont[3007] = 1'd0;
    assign memfont[3008] = 1'd0;
    assign memfont[3009] = 1'd0;
    assign memfont[3010] = 1'd0;
    assign memfont[3011] = 1'd0;
    assign memfont[3012] = 1'd0;
    assign memfont[3013] = 1'd0;
    assign memfont[3014] = 1'd0;
    assign memfont[3015] = 1'd0;
    assign memfont[3016] = 1'd0;
    assign memfont[3017] = 1'd1;
    assign memfont[3018] = 1'd1;
    assign memfont[3019] = 1'd0;
    assign memfont[3020] = 1'd0;
    assign memfont[3021] = 1'd0;
    assign memfont[3022] = 1'd0;
    assign memfont[3023] = 1'd0;
    assign memfont[3024] = 1'd0;
    assign memfont[3025] = 1'd1;
    assign memfont[3026] = 1'd1;
    assign memfont[3027] = 1'd0;
    assign memfont[3028] = 1'd0;
    assign memfont[3029] = 1'd0;
    assign memfont[3030] = 1'd0;
    assign memfont[3031] = 1'd0;
    assign memfont[3032] = 1'd0;
    assign memfont[3033] = 1'd1;
    assign memfont[3034] = 1'd1;
    assign memfont[3035] = 1'd0;
    assign memfont[3036] = 1'd0;
    assign memfont[3037] = 1'd0;
    assign memfont[3038] = 1'd1;
    assign memfont[3039] = 1'd1;
    assign memfont[3040] = 1'd0;
    assign memfont[3041] = 1'd0;
    assign memfont[3042] = 1'd0;
    assign memfont[3043] = 1'd1;
    assign memfont[3044] = 1'd1;
    assign memfont[3045] = 1'd0;
    assign memfont[3046] = 1'd0;
    assign memfont[3047] = 1'd0;
    assign memfont[3048] = 1'd0;
    assign memfont[3049] = 1'd1;
    assign memfont[3050] = 1'd1;
    assign memfont[3051] = 1'd0;
    assign memfont[3052] = 1'd1;
    assign memfont[3053] = 1'd0;
    assign memfont[3054] = 1'd1;
    assign memfont[3055] = 1'd1;
    assign memfont[3056] = 1'd0;
    assign memfont[3057] = 1'd1;
    assign memfont[3058] = 1'd1;
    assign memfont[3059] = 1'd0;
    assign memfont[3060] = 1'd0;
    assign memfont[3061] = 1'd0;
    assign memfont[3062] = 1'd0;
    assign memfont[3063] = 1'd0;
    assign memfont[3064] = 1'd1;
    assign memfont[3065] = 1'd1;
    assign memfont[3066] = 1'd1;
    assign memfont[3067] = 1'd0;
    assign memfont[3068] = 1'd0;
    assign memfont[3069] = 1'd0;
    assign memfont[3070] = 1'd0;
    assign memfont[3071] = 1'd0;
    assign memfont[3072] = 1'd0;
    assign memfont[3073] = 1'd0;
    assign memfont[3074] = 1'd0;
    assign memfont[3075] = 1'd0;
    assign memfont[3076] = 1'd1;
    assign memfont[3077] = 1'd1;
    assign memfont[3078] = 1'd1;
    assign memfont[3079] = 1'd1;
    assign memfont[3080] = 1'd0;
    assign memfont[3081] = 1'd0;
    assign memfont[3082] = 1'd0;
    assign memfont[3083] = 1'd0;
    assign memfont[3084] = 1'd0;
    assign memfont[3085] = 1'd0;
    assign memfont[3086] = 1'd0;
    assign memfont[3087] = 1'd0;
    assign memfont[3088] = 1'd0;
    assign memfont[3089] = 1'd1;
    assign memfont[3090] = 1'd1;
    assign memfont[3091] = 1'd0;
    assign memfont[3092] = 1'd0;
    assign memfont[3093] = 1'd0;
    assign memfont[3094] = 1'd0;
    assign memfont[3095] = 1'd0;
    assign memfont[3096] = 1'd0;
    assign memfont[3097] = 1'd0;
    assign memfont[3098] = 1'd0;
    assign memfont[3099] = 1'd0;
    assign memfont[3100] = 1'd0;
    assign memfont[3101] = 1'd1;
    assign memfont[3102] = 1'd1;
    assign memfont[3103] = 1'd0;
    assign memfont[3104] = 1'd0;
    assign memfont[3105] = 1'd0;
    assign memfont[3106] = 1'd0;
    assign memfont[3107] = 1'd0;
    assign memfont[3108] = 1'd0;
    assign memfont[3109] = 1'd1;
    assign memfont[3110] = 1'd1;
    assign memfont[3111] = 1'd0;
    assign memfont[3112] = 1'd0;
    assign memfont[3113] = 1'd1;
    assign memfont[3114] = 1'd1;
    assign memfont[3115] = 1'd0;
    assign memfont[3116] = 1'd0;
    assign memfont[3117] = 1'd1;
    assign memfont[3118] = 1'd1;
    assign memfont[3119] = 1'd0;
    assign memfont[3120] = 1'd0;
    assign memfont[3121] = 1'd1;
    assign memfont[3122] = 1'd1;
    assign memfont[3123] = 1'd0;
    assign memfont[3124] = 1'd0;
    assign memfont[3125] = 1'd0;
    assign memfont[3126] = 1'd0;
    assign memfont[3127] = 1'd0;
    assign memfont[3128] = 1'd0;
    assign memfont[3129] = 1'd1;
    assign memfont[3130] = 1'd1;
    assign memfont[3131] = 1'd0;
    assign memfont[3132] = 1'd0;
    assign memfont[3133] = 1'd0;
    assign memfont[3134] = 1'd0;
    assign memfont[3135] = 1'd1;
    assign memfont[3136] = 1'd1;
    assign memfont[3137] = 1'd0;
    assign memfont[3138] = 1'd0;
    assign memfont[3139] = 1'd1;
    assign memfont[3140] = 1'd1;
    assign memfont[3141] = 1'd0;
    assign memfont[3142] = 1'd0;
    assign memfont[3143] = 1'd0;
    assign memfont[3144] = 1'd0;
    assign memfont[3145] = 1'd1;
    assign memfont[3146] = 1'd1;
    assign memfont[3147] = 1'd1;
    assign memfont[3148] = 1'd1;
    assign memfont[3149] = 1'd1;
    assign memfont[3150] = 1'd1;
    assign memfont[3151] = 1'd1;
    assign memfont[3152] = 1'd1;
    assign memfont[3153] = 1'd0;
    assign memfont[3154] = 1'd0;
    assign memfont[3155] = 1'd0;
    assign memfont[3156] = 1'd0;
    assign memfont[3157] = 1'd1;
    assign memfont[3158] = 1'd1;
    assign memfont[3159] = 1'd0;
    assign memfont[3160] = 1'd0;
    assign memfont[3161] = 1'd0;
    assign memfont[3162] = 1'd0;
    assign memfont[3163] = 1'd0;
    assign memfont[3164] = 1'd0;
    assign memfont[3165] = 1'd0;
    assign memfont[3166] = 1'd0;
    assign memfont[3167] = 1'd0;
    assign memfont[3168] = 1'd0;
    assign memfont[3169] = 1'd1;
    assign memfont[3170] = 1'd1;
    assign memfont[3171] = 1'd0;
    assign memfont[3172] = 1'd0;
    assign memfont[3173] = 1'd0;
    assign memfont[3174] = 1'd0;
    assign memfont[3175] = 1'd0;
    assign memfont[3176] = 1'd0;
    assign memfont[3177] = 1'd1;
    assign memfont[3178] = 1'd1;
    assign memfont[3179] = 1'd0;
    assign memfont[3180] = 1'd0;
    assign memfont[3181] = 1'd1;
    assign memfont[3182] = 1'd1;
    assign memfont[3183] = 1'd1;
    assign memfont[3184] = 1'd1;
    assign memfont[3185] = 1'd1;
    assign memfont[3186] = 1'd1;
    assign memfont[3187] = 1'd1;
    assign memfont[3188] = 1'd1;
    assign memfont[3189] = 1'd1;
    assign memfont[3190] = 1'd0;
    assign memfont[3191] = 1'd0;
    assign memfont[3192] = 1'd0;
    assign memfont[3193] = 1'd1;
    assign memfont[3194] = 1'd1;
    assign memfont[3195] = 1'd1;
    assign memfont[3196] = 1'd1;
    assign memfont[3197] = 1'd1;
    assign memfont[3198] = 1'd1;
    assign memfont[3199] = 1'd1;
    assign memfont[3200] = 1'd1;
    assign memfont[3201] = 1'd0;
    assign memfont[3202] = 1'd0;
    assign memfont[3203] = 1'd0;
    assign memfont[3204] = 1'd0;
    assign memfont[3205] = 1'd1;
    assign memfont[3206] = 1'd1;
    assign memfont[3207] = 1'd0;
    assign memfont[3208] = 1'd0;
    assign memfont[3209] = 1'd0;
    assign memfont[3210] = 1'd1;
    assign memfont[3211] = 1'd1;
    assign memfont[3212] = 1'd1;
    assign memfont[3213] = 1'd1;
    assign memfont[3214] = 1'd1;
    assign memfont[3215] = 1'd0;
    assign memfont[3216] = 1'd0;
    assign memfont[3217] = 1'd1;
    assign memfont[3218] = 1'd1;
    assign memfont[3219] = 1'd1;
    assign memfont[3220] = 1'd1;
    assign memfont[3221] = 1'd1;
    assign memfont[3222] = 1'd1;
    assign memfont[3223] = 1'd1;
    assign memfont[3224] = 1'd1;
    assign memfont[3225] = 1'd1;
    assign memfont[3226] = 1'd1;
    assign memfont[3227] = 1'd0;
    assign memfont[3228] = 1'd0;
    assign memfont[3229] = 1'd0;
    assign memfont[3230] = 1'd0;
    assign memfont[3231] = 1'd0;
    assign memfont[3232] = 1'd0;
    assign memfont[3233] = 1'd1;
    assign memfont[3234] = 1'd1;
    assign memfont[3235] = 1'd0;
    assign memfont[3236] = 1'd0;
    assign memfont[3237] = 1'd0;
    assign memfont[3238] = 1'd0;
    assign memfont[3239] = 1'd0;
    assign memfont[3240] = 1'd0;
    assign memfont[3241] = 1'd0;
    assign memfont[3242] = 1'd0;
    assign memfont[3243] = 1'd0;
    assign memfont[3244] = 1'd0;
    assign memfont[3245] = 1'd0;
    assign memfont[3246] = 1'd0;
    assign memfont[3247] = 1'd0;
    assign memfont[3248] = 1'd1;
    assign memfont[3249] = 1'd1;
    assign memfont[3250] = 1'd1;
    assign memfont[3251] = 1'd0;
    assign memfont[3252] = 1'd0;
    assign memfont[3253] = 1'd1;
    assign memfont[3254] = 1'd1;
    assign memfont[3255] = 1'd1;
    assign memfont[3256] = 1'd1;
    assign memfont[3257] = 1'd1;
    assign memfont[3258] = 1'd1;
    assign memfont[3259] = 1'd0;
    assign memfont[3260] = 1'd0;
    assign memfont[3261] = 1'd0;
    assign memfont[3262] = 1'd0;
    assign memfont[3263] = 1'd0;
    assign memfont[3264] = 1'd0;
    assign memfont[3265] = 1'd1;
    assign memfont[3266] = 1'd1;
    assign memfont[3267] = 1'd0;
    assign memfont[3268] = 1'd0;
    assign memfont[3269] = 1'd0;
    assign memfont[3270] = 1'd0;
    assign memfont[3271] = 1'd0;
    assign memfont[3272] = 1'd0;
    assign memfont[3273] = 1'd0;
    assign memfont[3274] = 1'd0;
    assign memfont[3275] = 1'd0;
    assign memfont[3276] = 1'd0;
    assign memfont[3277] = 1'd1;
    assign memfont[3278] = 1'd1;
    assign memfont[3279] = 1'd0;
    assign memfont[3280] = 1'd1;
    assign memfont[3281] = 1'd0;
    assign memfont[3282] = 1'd0;
    assign memfont[3283] = 1'd1;
    assign memfont[3284] = 1'd0;
    assign memfont[3285] = 1'd1;
    assign memfont[3286] = 1'd1;
    assign memfont[3287] = 1'd0;
    assign memfont[3288] = 1'd0;
    assign memfont[3289] = 1'd1;
    assign memfont[3290] = 1'd1;
    assign memfont[3291] = 1'd0;
    assign memfont[3292] = 1'd0;
    assign memfont[3293] = 1'd1;
    assign memfont[3294] = 1'd1;
    assign memfont[3295] = 1'd0;
    assign memfont[3296] = 1'd0;
    assign memfont[3297] = 1'd1;
    assign memfont[3298] = 1'd1;
    assign memfont[3299] = 1'd0;
    assign memfont[3300] = 1'd0;
    assign memfont[3301] = 1'd1;
    assign memfont[3302] = 1'd1;
    assign memfont[3303] = 1'd0;
    assign memfont[3304] = 1'd0;
    assign memfont[3305] = 1'd0;
    assign memfont[3306] = 1'd0;
    assign memfont[3307] = 1'd0;
    assign memfont[3308] = 1'd0;
    assign memfont[3309] = 1'd1;
    assign memfont[3310] = 1'd1;
    assign memfont[3311] = 1'd0;
    assign memfont[3312] = 1'd0;
    assign memfont[3313] = 1'd1;
    assign memfont[3314] = 1'd1;
    assign memfont[3315] = 1'd1;
    assign memfont[3316] = 1'd1;
    assign memfont[3317] = 1'd1;
    assign memfont[3318] = 1'd1;
    assign memfont[3319] = 1'd1;
    assign memfont[3320] = 1'd1;
    assign memfont[3321] = 1'd1;
    assign memfont[3322] = 1'd0;
    assign memfont[3323] = 1'd0;
    assign memfont[3324] = 1'd0;
    assign memfont[3325] = 1'd1;
    assign memfont[3326] = 1'd1;
    assign memfont[3327] = 1'd0;
    assign memfont[3328] = 1'd0;
    assign memfont[3329] = 1'd0;
    assign memfont[3330] = 1'd0;
    assign memfont[3331] = 1'd0;
    assign memfont[3332] = 1'd0;
    assign memfont[3333] = 1'd1;
    assign memfont[3334] = 1'd1;
    assign memfont[3335] = 1'd0;
    assign memfont[3336] = 1'd0;
    assign memfont[3337] = 1'd1;
    assign memfont[3338] = 1'd1;
    assign memfont[3339] = 1'd1;
    assign memfont[3340] = 1'd1;
    assign memfont[3341] = 1'd1;
    assign memfont[3342] = 1'd1;
    assign memfont[3343] = 1'd1;
    assign memfont[3344] = 1'd1;
    assign memfont[3345] = 1'd0;
    assign memfont[3346] = 1'd0;
    assign memfont[3347] = 1'd0;
    assign memfont[3348] = 1'd0;
    assign memfont[3349] = 1'd0;
    assign memfont[3350] = 1'd0;
    assign memfont[3351] = 1'd0;
    assign memfont[3352] = 1'd1;
    assign memfont[3353] = 1'd1;
    assign memfont[3354] = 1'd1;
    assign memfont[3355] = 1'd1;
    assign memfont[3356] = 1'd1;
    assign memfont[3357] = 1'd0;
    assign memfont[3358] = 1'd0;
    assign memfont[3359] = 1'd0;
    assign memfont[3360] = 1'd0;
    assign memfont[3361] = 1'd0;
    assign memfont[3362] = 1'd0;
    assign memfont[3363] = 1'd0;
    assign memfont[3364] = 1'd0;
    assign memfont[3365] = 1'd1;
    assign memfont[3366] = 1'd1;
    assign memfont[3367] = 1'd0;
    assign memfont[3368] = 1'd0;
    assign memfont[3369] = 1'd0;
    assign memfont[3370] = 1'd0;
    assign memfont[3371] = 1'd0;
    assign memfont[3372] = 1'd0;
    assign memfont[3373] = 1'd1;
    assign memfont[3374] = 1'd1;
    assign memfont[3375] = 1'd0;
    assign memfont[3376] = 1'd0;
    assign memfont[3377] = 1'd0;
    assign memfont[3378] = 1'd0;
    assign memfont[3379] = 1'd0;
    assign memfont[3380] = 1'd0;
    assign memfont[3381] = 1'd1;
    assign memfont[3382] = 1'd1;
    assign memfont[3383] = 1'd0;
    assign memfont[3384] = 1'd0;
    assign memfont[3385] = 1'd0;
    assign memfont[3386] = 1'd1;
    assign memfont[3387] = 1'd1;
    assign memfont[3388] = 1'd1;
    assign memfont[3389] = 1'd0;
    assign memfont[3390] = 1'd0;
    assign memfont[3391] = 1'd1;
    assign memfont[3392] = 1'd1;
    assign memfont[3393] = 1'd0;
    assign memfont[3394] = 1'd0;
    assign memfont[3395] = 1'd0;
    assign memfont[3396] = 1'd0;
    assign memfont[3397] = 1'd1;
    assign memfont[3398] = 1'd1;
    assign memfont[3399] = 1'd0;
    assign memfont[3400] = 1'd1;
    assign memfont[3401] = 1'd0;
    assign memfont[3402] = 1'd1;
    assign memfont[3403] = 1'd1;
    assign memfont[3404] = 1'd0;
    assign memfont[3405] = 1'd1;
    assign memfont[3406] = 1'd1;
    assign memfont[3407] = 1'd0;
    assign memfont[3408] = 1'd0;
    assign memfont[3409] = 1'd0;
    assign memfont[3410] = 1'd0;
    assign memfont[3411] = 1'd0;
    assign memfont[3412] = 1'd0;
    assign memfont[3413] = 1'd1;
    assign memfont[3414] = 1'd1;
    assign memfont[3415] = 1'd0;
    assign memfont[3416] = 1'd0;
    assign memfont[3417] = 1'd0;
    assign memfont[3418] = 1'd0;
    assign memfont[3419] = 1'd0;
    assign memfont[3420] = 1'd0;
    assign memfont[3421] = 1'd0;
    assign memfont[3422] = 1'd0;
    assign memfont[3423] = 1'd0;
    assign memfont[3424] = 1'd1;
    assign memfont[3425] = 1'd1;
    assign memfont[3426] = 1'd1;
    assign memfont[3427] = 1'd0;
    assign memfont[3428] = 1'd0;
    assign memfont[3429] = 1'd0;
    assign memfont[3430] = 1'd0;
    assign memfont[3431] = 1'd0;
    assign memfont[3432] = 1'd0;
    assign memfont[3433] = 1'd0;
    assign memfont[3434] = 1'd0;
    assign memfont[3435] = 1'd0;
    assign memfont[3436] = 1'd0;
    assign memfont[3437] = 1'd1;
    assign memfont[3438] = 1'd1;
    assign memfont[3439] = 1'd0;
    assign memfont[3440] = 1'd0;
    assign memfont[3441] = 1'd0;
    assign memfont[3442] = 1'd0;
    assign memfont[3443] = 1'd0;
    assign memfont[3444] = 1'd0;
    assign memfont[3445] = 1'd0;
    assign memfont[3446] = 1'd0;
    assign memfont[3447] = 1'd0;
    assign memfont[3448] = 1'd0;
    assign memfont[3449] = 1'd1;
    assign memfont[3450] = 1'd1;
    assign memfont[3451] = 1'd0;
    assign memfont[3452] = 1'd0;
    assign memfont[3453] = 1'd0;
    assign memfont[3454] = 1'd0;
    assign memfont[3455] = 1'd0;
    assign memfont[3456] = 1'd0;
    assign memfont[3457] = 1'd1;
    assign memfont[3458] = 1'd1;
    assign memfont[3459] = 1'd1;
    assign memfont[3460] = 1'd1;
    assign memfont[3461] = 1'd1;
    assign memfont[3462] = 1'd1;
    assign memfont[3463] = 1'd0;
    assign memfont[3464] = 1'd0;
    assign memfont[3465] = 1'd1;
    assign memfont[3466] = 1'd1;
    assign memfont[3467] = 1'd0;
    assign memfont[3468] = 1'd0;
    assign memfont[3469] = 1'd1;
    assign memfont[3470] = 1'd1;
    assign memfont[3471] = 1'd1;
    assign memfont[3472] = 1'd1;
    assign memfont[3473] = 1'd0;
    assign memfont[3474] = 1'd0;
    assign memfont[3475] = 1'd1;
    assign memfont[3476] = 1'd1;
    assign memfont[3477] = 1'd1;
    assign memfont[3478] = 1'd1;
    assign memfont[3479] = 1'd0;
    assign memfont[3480] = 1'd0;
    assign memfont[3481] = 1'd0;
    assign memfont[3482] = 1'd1;
    assign memfont[3483] = 1'd1;
    assign memfont[3484] = 1'd0;
    assign memfont[3485] = 1'd0;
    assign memfont[3486] = 1'd0;
    assign memfont[3487] = 1'd1;
    assign memfont[3488] = 1'd1;
    assign memfont[3489] = 1'd0;
    assign memfont[3490] = 1'd0;
    assign memfont[3491] = 1'd0;
    assign memfont[3492] = 1'd0;
    assign memfont[3493] = 1'd1;
    assign memfont[3494] = 1'd1;
    assign memfont[3495] = 1'd0;
    assign memfont[3496] = 1'd0;
    assign memfont[3497] = 1'd0;
    assign memfont[3498] = 1'd0;
    assign memfont[3499] = 1'd0;
    assign memfont[3500] = 1'd1;
    assign memfont[3501] = 1'd1;
    assign memfont[3502] = 1'd0;
    assign memfont[3503] = 1'd0;
    assign memfont[3504] = 1'd0;
    assign memfont[3505] = 1'd1;
    assign memfont[3506] = 1'd1;
    assign memfont[3507] = 1'd0;
    assign memfont[3508] = 1'd0;
    assign memfont[3509] = 1'd0;
    assign memfont[3510] = 1'd0;
    assign memfont[3511] = 1'd0;
    assign memfont[3512] = 1'd0;
    assign memfont[3513] = 1'd0;
    assign memfont[3514] = 1'd0;
    assign memfont[3515] = 1'd0;
    assign memfont[3516] = 1'd0;
    assign memfont[3517] = 1'd1;
    assign memfont[3518] = 1'd1;
    assign memfont[3519] = 1'd0;
    assign memfont[3520] = 1'd0;
    assign memfont[3521] = 1'd0;
    assign memfont[3522] = 1'd0;
    assign memfont[3523] = 1'd0;
    assign memfont[3524] = 1'd0;
    assign memfont[3525] = 1'd1;
    assign memfont[3526] = 1'd1;
    assign memfont[3527] = 1'd0;
    assign memfont[3528] = 1'd0;
    assign memfont[3529] = 1'd1;
    assign memfont[3530] = 1'd1;
    assign memfont[3531] = 1'd0;
    assign memfont[3532] = 1'd0;
    assign memfont[3533] = 1'd0;
    assign memfont[3534] = 1'd0;
    assign memfont[3535] = 1'd0;
    assign memfont[3536] = 1'd0;
    assign memfont[3537] = 1'd0;
    assign memfont[3538] = 1'd0;
    assign memfont[3539] = 1'd0;
    assign memfont[3540] = 1'd0;
    assign memfont[3541] = 1'd1;
    assign memfont[3542] = 1'd1;
    assign memfont[3543] = 1'd0;
    assign memfont[3544] = 1'd0;
    assign memfont[3545] = 1'd0;
    assign memfont[3546] = 1'd0;
    assign memfont[3547] = 1'd0;
    assign memfont[3548] = 1'd0;
    assign memfont[3549] = 1'd0;
    assign memfont[3550] = 1'd0;
    assign memfont[3551] = 1'd0;
    assign memfont[3552] = 1'd0;
    assign memfont[3553] = 1'd1;
    assign memfont[3554] = 1'd1;
    assign memfont[3555] = 1'd0;
    assign memfont[3556] = 1'd0;
    assign memfont[3557] = 1'd0;
    assign memfont[3558] = 1'd1;
    assign memfont[3559] = 1'd1;
    assign memfont[3560] = 1'd1;
    assign memfont[3561] = 1'd1;
    assign memfont[3562] = 1'd1;
    assign memfont[3563] = 1'd0;
    assign memfont[3564] = 1'd0;
    assign memfont[3565] = 1'd1;
    assign memfont[3566] = 1'd1;
    assign memfont[3567] = 1'd0;
    assign memfont[3568] = 1'd0;
    assign memfont[3569] = 1'd0;
    assign memfont[3570] = 1'd0;
    assign memfont[3571] = 1'd0;
    assign memfont[3572] = 1'd0;
    assign memfont[3573] = 1'd1;
    assign memfont[3574] = 1'd1;
    assign memfont[3575] = 1'd0;
    assign memfont[3576] = 1'd0;
    assign memfont[3577] = 1'd0;
    assign memfont[3578] = 1'd0;
    assign memfont[3579] = 1'd0;
    assign memfont[3580] = 1'd0;
    assign memfont[3581] = 1'd1;
    assign memfont[3582] = 1'd1;
    assign memfont[3583] = 1'd0;
    assign memfont[3584] = 1'd0;
    assign memfont[3585] = 1'd0;
    assign memfont[3586] = 1'd0;
    assign memfont[3587] = 1'd0;
    assign memfont[3588] = 1'd0;
    assign memfont[3589] = 1'd0;
    assign memfont[3590] = 1'd0;
    assign memfont[3591] = 1'd0;
    assign memfont[3592] = 1'd0;
    assign memfont[3593] = 1'd0;
    assign memfont[3594] = 1'd0;
    assign memfont[3595] = 1'd0;
    assign memfont[3596] = 1'd1;
    assign memfont[3597] = 1'd1;
    assign memfont[3598] = 1'd1;
    assign memfont[3599] = 1'd0;
    assign memfont[3600] = 1'd0;
    assign memfont[3601] = 1'd1;
    assign memfont[3602] = 1'd1;
    assign memfont[3603] = 1'd1;
    assign memfont[3604] = 1'd0;
    assign memfont[3605] = 1'd1;
    assign memfont[3606] = 1'd1;
    assign memfont[3607] = 1'd1;
    assign memfont[3608] = 1'd0;
    assign memfont[3609] = 1'd0;
    assign memfont[3610] = 1'd0;
    assign memfont[3611] = 1'd0;
    assign memfont[3612] = 1'd0;
    assign memfont[3613] = 1'd1;
    assign memfont[3614] = 1'd1;
    assign memfont[3615] = 1'd0;
    assign memfont[3616] = 1'd0;
    assign memfont[3617] = 1'd0;
    assign memfont[3618] = 1'd0;
    assign memfont[3619] = 1'd0;
    assign memfont[3620] = 1'd0;
    assign memfont[3621] = 1'd0;
    assign memfont[3622] = 1'd0;
    assign memfont[3623] = 1'd0;
    assign memfont[3624] = 1'd0;
    assign memfont[3625] = 1'd1;
    assign memfont[3626] = 1'd1;
    assign memfont[3627] = 1'd0;
    assign memfont[3628] = 1'd1;
    assign memfont[3629] = 1'd1;
    assign memfont[3630] = 1'd1;
    assign memfont[3631] = 1'd1;
    assign memfont[3632] = 1'd0;
    assign memfont[3633] = 1'd1;
    assign memfont[3634] = 1'd1;
    assign memfont[3635] = 1'd0;
    assign memfont[3636] = 1'd0;
    assign memfont[3637] = 1'd1;
    assign memfont[3638] = 1'd1;
    assign memfont[3639] = 1'd0;
    assign memfont[3640] = 1'd0;
    assign memfont[3641] = 1'd1;
    assign memfont[3642] = 1'd1;
    assign memfont[3643] = 1'd0;
    assign memfont[3644] = 1'd0;
    assign memfont[3645] = 1'd1;
    assign memfont[3646] = 1'd1;
    assign memfont[3647] = 1'd0;
    assign memfont[3648] = 1'd0;
    assign memfont[3649] = 1'd1;
    assign memfont[3650] = 1'd1;
    assign memfont[3651] = 1'd0;
    assign memfont[3652] = 1'd0;
    assign memfont[3653] = 1'd0;
    assign memfont[3654] = 1'd0;
    assign memfont[3655] = 1'd0;
    assign memfont[3656] = 1'd0;
    assign memfont[3657] = 1'd1;
    assign memfont[3658] = 1'd1;
    assign memfont[3659] = 1'd0;
    assign memfont[3660] = 1'd0;
    assign memfont[3661] = 1'd1;
    assign memfont[3662] = 1'd1;
    assign memfont[3663] = 1'd1;
    assign memfont[3664] = 1'd1;
    assign memfont[3665] = 1'd1;
    assign memfont[3666] = 1'd1;
    assign memfont[3667] = 1'd1;
    assign memfont[3668] = 1'd1;
    assign memfont[3669] = 1'd0;
    assign memfont[3670] = 1'd0;
    assign memfont[3671] = 1'd0;
    assign memfont[3672] = 1'd0;
    assign memfont[3673] = 1'd1;
    assign memfont[3674] = 1'd1;
    assign memfont[3675] = 1'd0;
    assign memfont[3676] = 1'd0;
    assign memfont[3677] = 1'd0;
    assign memfont[3678] = 1'd0;
    assign memfont[3679] = 1'd0;
    assign memfont[3680] = 1'd0;
    assign memfont[3681] = 1'd1;
    assign memfont[3682] = 1'd1;
    assign memfont[3683] = 1'd0;
    assign memfont[3684] = 1'd0;
    assign memfont[3685] = 1'd1;
    assign memfont[3686] = 1'd1;
    assign memfont[3687] = 1'd1;
    assign memfont[3688] = 1'd1;
    assign memfont[3689] = 1'd1;
    assign memfont[3690] = 1'd1;
    assign memfont[3691] = 1'd1;
    assign memfont[3692] = 1'd0;
    assign memfont[3693] = 1'd0;
    assign memfont[3694] = 1'd0;
    assign memfont[3695] = 1'd0;
    assign memfont[3696] = 1'd0;
    assign memfont[3697] = 1'd0;
    assign memfont[3698] = 1'd0;
    assign memfont[3699] = 1'd0;
    assign memfont[3700] = 1'd0;
    assign memfont[3701] = 1'd0;
    assign memfont[3702] = 1'd1;
    assign memfont[3703] = 1'd1;
    assign memfont[3704] = 1'd1;
    assign memfont[3705] = 1'd1;
    assign memfont[3706] = 1'd0;
    assign memfont[3707] = 1'd0;
    assign memfont[3708] = 1'd0;
    assign memfont[3709] = 1'd0;
    assign memfont[3710] = 1'd0;
    assign memfont[3711] = 1'd0;
    assign memfont[3712] = 1'd0;
    assign memfont[3713] = 1'd1;
    assign memfont[3714] = 1'd1;
    assign memfont[3715] = 1'd0;
    assign memfont[3716] = 1'd0;
    assign memfont[3717] = 1'd0;
    assign memfont[3718] = 1'd0;
    assign memfont[3719] = 1'd0;
    assign memfont[3720] = 1'd0;
    assign memfont[3721] = 1'd1;
    assign memfont[3722] = 1'd1;
    assign memfont[3723] = 1'd0;
    assign memfont[3724] = 1'd0;
    assign memfont[3725] = 1'd0;
    assign memfont[3726] = 1'd0;
    assign memfont[3727] = 1'd0;
    assign memfont[3728] = 1'd0;
    assign memfont[3729] = 1'd1;
    assign memfont[3730] = 1'd1;
    assign memfont[3731] = 1'd0;
    assign memfont[3732] = 1'd0;
    assign memfont[3733] = 1'd0;
    assign memfont[3734] = 1'd0;
    assign memfont[3735] = 1'd1;
    assign memfont[3736] = 1'd1;
    assign memfont[3737] = 1'd0;
    assign memfont[3738] = 1'd0;
    assign memfont[3739] = 1'd1;
    assign memfont[3740] = 1'd1;
    assign memfont[3741] = 1'd0;
    assign memfont[3742] = 1'd0;
    assign memfont[3743] = 1'd0;
    assign memfont[3744] = 1'd0;
    assign memfont[3745] = 1'd1;
    assign memfont[3746] = 1'd1;
    assign memfont[3747] = 1'd0;
    assign memfont[3748] = 1'd1;
    assign memfont[3749] = 1'd0;
    assign memfont[3750] = 1'd0;
    assign memfont[3751] = 1'd1;
    assign memfont[3752] = 1'd0;
    assign memfont[3753] = 1'd1;
    assign memfont[3754] = 1'd0;
    assign memfont[3755] = 1'd0;
    assign memfont[3756] = 1'd0;
    assign memfont[3757] = 1'd0;
    assign memfont[3758] = 1'd0;
    assign memfont[3759] = 1'd0;
    assign memfont[3760] = 1'd1;
    assign memfont[3761] = 1'd1;
    assign memfont[3762] = 1'd1;
    assign memfont[3763] = 1'd1;
    assign memfont[3764] = 1'd0;
    assign memfont[3765] = 1'd0;
    assign memfont[3766] = 1'd0;
    assign memfont[3767] = 1'd0;
    assign memfont[3768] = 1'd0;
    assign memfont[3769] = 1'd0;
    assign memfont[3770] = 1'd0;
    assign memfont[3771] = 1'd0;
    assign memfont[3772] = 1'd0;
    assign memfont[3773] = 1'd1;
    assign memfont[3774] = 1'd1;
    assign memfont[3775] = 1'd0;
    assign memfont[3776] = 1'd0;
    assign memfont[3777] = 1'd0;
    assign memfont[3778] = 1'd0;
    assign memfont[3779] = 1'd0;
    assign memfont[3780] = 1'd0;
    assign memfont[3781] = 1'd0;
    assign memfont[3782] = 1'd0;
    assign memfont[3783] = 1'd0;
    assign memfont[3784] = 1'd1;
    assign memfont[3785] = 1'd1;
    assign memfont[3786] = 1'd0;
    assign memfont[3787] = 1'd0;
    assign memfont[3788] = 1'd0;
    assign memfont[3789] = 1'd0;
    assign memfont[3790] = 1'd0;
    assign memfont[3791] = 1'd0;
    assign memfont[3792] = 1'd0;
    assign memfont[3793] = 1'd0;
    assign memfont[3794] = 1'd0;
    assign memfont[3795] = 1'd0;
    assign memfont[3796] = 1'd0;
    assign memfont[3797] = 1'd1;
    assign memfont[3798] = 1'd1;
    assign memfont[3799] = 1'd0;
    assign memfont[3800] = 1'd0;
    assign memfont[3801] = 1'd0;
    assign memfont[3802] = 1'd0;
    assign memfont[3803] = 1'd0;
    assign memfont[3804] = 1'd0;
    assign memfont[3805] = 1'd1;
    assign memfont[3806] = 1'd1;
    assign memfont[3807] = 1'd0;
    assign memfont[3808] = 1'd0;
    assign memfont[3809] = 1'd1;
    assign memfont[3810] = 1'd1;
    assign memfont[3811] = 1'd0;
    assign memfont[3812] = 1'd0;
    assign memfont[3813] = 1'd1;
    assign memfont[3814] = 1'd1;
    assign memfont[3815] = 1'd0;
    assign memfont[3816] = 1'd0;
    assign memfont[3817] = 1'd1;
    assign memfont[3818] = 1'd1;
    assign memfont[3819] = 1'd1;
    assign memfont[3820] = 1'd1;
    assign memfont[3821] = 1'd0;
    assign memfont[3822] = 1'd0;
    assign memfont[3823] = 1'd1;
    assign memfont[3824] = 1'd1;
    assign memfont[3825] = 1'd1;
    assign memfont[3826] = 1'd1;
    assign memfont[3827] = 1'd0;
    assign memfont[3828] = 1'd0;
    assign memfont[3829] = 1'd0;
    assign memfont[3830] = 1'd1;
    assign memfont[3831] = 1'd1;
    assign memfont[3832] = 1'd1;
    assign memfont[3833] = 1'd1;
    assign memfont[3834] = 1'd1;
    assign memfont[3835] = 1'd1;
    assign memfont[3836] = 1'd1;
    assign memfont[3837] = 1'd1;
    assign memfont[3838] = 1'd0;
    assign memfont[3839] = 1'd0;
    assign memfont[3840] = 1'd0;
    assign memfont[3841] = 1'd1;
    assign memfont[3842] = 1'd1;
    assign memfont[3843] = 1'd0;
    assign memfont[3844] = 1'd0;
    assign memfont[3845] = 1'd0;
    assign memfont[3846] = 1'd0;
    assign memfont[3847] = 1'd0;
    assign memfont[3848] = 1'd0;
    assign memfont[3849] = 1'd1;
    assign memfont[3850] = 1'd1;
    assign memfont[3851] = 1'd0;
    assign memfont[3852] = 1'd0;
    assign memfont[3853] = 1'd1;
    assign memfont[3854] = 1'd1;
    assign memfont[3855] = 1'd0;
    assign memfont[3856] = 1'd0;
    assign memfont[3857] = 1'd0;
    assign memfont[3858] = 1'd0;
    assign memfont[3859] = 1'd0;
    assign memfont[3860] = 1'd0;
    assign memfont[3861] = 1'd1;
    assign memfont[3862] = 1'd1;
    assign memfont[3863] = 1'd0;
    assign memfont[3864] = 1'd0;
    assign memfont[3865] = 1'd1;
    assign memfont[3866] = 1'd1;
    assign memfont[3867] = 1'd0;
    assign memfont[3868] = 1'd0;
    assign memfont[3869] = 1'd0;
    assign memfont[3870] = 1'd0;
    assign memfont[3871] = 1'd0;
    assign memfont[3872] = 1'd0;
    assign memfont[3873] = 1'd1;
    assign memfont[3874] = 1'd1;
    assign memfont[3875] = 1'd0;
    assign memfont[3876] = 1'd0;
    assign memfont[3877] = 1'd1;
    assign memfont[3878] = 1'd1;
    assign memfont[3879] = 1'd0;
    assign memfont[3880] = 1'd0;
    assign memfont[3881] = 1'd0;
    assign memfont[3882] = 1'd0;
    assign memfont[3883] = 1'd0;
    assign memfont[3884] = 1'd0;
    assign memfont[3885] = 1'd0;
    assign memfont[3886] = 1'd0;
    assign memfont[3887] = 1'd0;
    assign memfont[3888] = 1'd0;
    assign memfont[3889] = 1'd1;
    assign memfont[3890] = 1'd1;
    assign memfont[3891] = 1'd0;
    assign memfont[3892] = 1'd0;
    assign memfont[3893] = 1'd0;
    assign memfont[3894] = 1'd0;
    assign memfont[3895] = 1'd0;
    assign memfont[3896] = 1'd0;
    assign memfont[3897] = 1'd0;
    assign memfont[3898] = 1'd0;
    assign memfont[3899] = 1'd0;
    assign memfont[3900] = 1'd0;
    assign memfont[3901] = 1'd1;
    assign memfont[3902] = 1'd1;
    assign memfont[3903] = 1'd0;
    assign memfont[3904] = 1'd0;
    assign memfont[3905] = 1'd0;
    assign memfont[3906] = 1'd0;
    assign memfont[3907] = 1'd0;
    assign memfont[3908] = 1'd0;
    assign memfont[3909] = 1'd1;
    assign memfont[3910] = 1'd1;
    assign memfont[3911] = 1'd0;
    assign memfont[3912] = 1'd0;
    assign memfont[3913] = 1'd1;
    assign memfont[3914] = 1'd1;
    assign memfont[3915] = 1'd0;
    assign memfont[3916] = 1'd0;
    assign memfont[3917] = 1'd0;
    assign memfont[3918] = 1'd0;
    assign memfont[3919] = 1'd0;
    assign memfont[3920] = 1'd0;
    assign memfont[3921] = 1'd1;
    assign memfont[3922] = 1'd1;
    assign memfont[3923] = 1'd0;
    assign memfont[3924] = 1'd0;
    assign memfont[3925] = 1'd0;
    assign memfont[3926] = 1'd0;
    assign memfont[3927] = 1'd0;
    assign memfont[3928] = 1'd0;
    assign memfont[3929] = 1'd1;
    assign memfont[3930] = 1'd1;
    assign memfont[3931] = 1'd0;
    assign memfont[3932] = 1'd0;
    assign memfont[3933] = 1'd0;
    assign memfont[3934] = 1'd0;
    assign memfont[3935] = 1'd0;
    assign memfont[3936] = 1'd0;
    assign memfont[3937] = 1'd1;
    assign memfont[3938] = 1'd1;
    assign memfont[3939] = 1'd0;
    assign memfont[3940] = 1'd0;
    assign memfont[3941] = 1'd0;
    assign memfont[3942] = 1'd0;
    assign memfont[3943] = 1'd0;
    assign memfont[3944] = 1'd1;
    assign memfont[3945] = 1'd1;
    assign memfont[3946] = 1'd1;
    assign memfont[3947] = 1'd0;
    assign memfont[3948] = 1'd0;
    assign memfont[3949] = 1'd1;
    assign memfont[3950] = 1'd1;
    assign memfont[3951] = 1'd0;
    assign memfont[3952] = 1'd0;
    assign memfont[3953] = 1'd0;
    assign memfont[3954] = 1'd1;
    assign memfont[3955] = 1'd1;
    assign memfont[3956] = 1'd0;
    assign memfont[3957] = 1'd0;
    assign memfont[3958] = 1'd0;
    assign memfont[3959] = 1'd0;
    assign memfont[3960] = 1'd0;
    assign memfont[3961] = 1'd1;
    assign memfont[3962] = 1'd1;
    assign memfont[3963] = 1'd0;
    assign memfont[3964] = 1'd0;
    assign memfont[3965] = 1'd0;
    assign memfont[3966] = 1'd0;
    assign memfont[3967] = 1'd0;
    assign memfont[3968] = 1'd0;
    assign memfont[3969] = 1'd0;
    assign memfont[3970] = 1'd0;
    assign memfont[3971] = 1'd0;
    assign memfont[3972] = 1'd0;
    assign memfont[3973] = 1'd1;
    assign memfont[3974] = 1'd1;
    assign memfont[3975] = 1'd0;
    assign memfont[3976] = 1'd1;
    assign memfont[3977] = 1'd1;
    assign memfont[3978] = 1'd1;
    assign memfont[3979] = 1'd1;
    assign memfont[3980] = 1'd0;
    assign memfont[3981] = 1'd1;
    assign memfont[3982] = 1'd1;
    assign memfont[3983] = 1'd0;
    assign memfont[3984] = 1'd0;
    assign memfont[3985] = 1'd1;
    assign memfont[3986] = 1'd1;
    assign memfont[3987] = 1'd0;
    assign memfont[3988] = 1'd0;
    assign memfont[3989] = 1'd0;
    assign memfont[3990] = 1'd1;
    assign memfont[3991] = 1'd1;
    assign memfont[3992] = 1'd0;
    assign memfont[3993] = 1'd1;
    assign memfont[3994] = 1'd1;
    assign memfont[3995] = 1'd0;
    assign memfont[3996] = 1'd0;
    assign memfont[3997] = 1'd1;
    assign memfont[3998] = 1'd1;
    assign memfont[3999] = 1'd0;
    assign memfont[4000] = 1'd0;
    assign memfont[4001] = 1'd0;
    assign memfont[4002] = 1'd0;
    assign memfont[4003] = 1'd0;
    assign memfont[4004] = 1'd0;
    assign memfont[4005] = 1'd1;
    assign memfont[4006] = 1'd1;
    assign memfont[4007] = 1'd0;
    assign memfont[4008] = 1'd0;
    assign memfont[4009] = 1'd1;
    assign memfont[4010] = 1'd1;
    assign memfont[4011] = 1'd0;
    assign memfont[4012] = 1'd0;
    assign memfont[4013] = 1'd0;
    assign memfont[4014] = 1'd0;
    assign memfont[4015] = 1'd0;
    assign memfont[4016] = 1'd0;
    assign memfont[4017] = 1'd0;
    assign memfont[4018] = 1'd0;
    assign memfont[4019] = 1'd0;
    assign memfont[4020] = 1'd0;
    assign memfont[4021] = 1'd1;
    assign memfont[4022] = 1'd1;
    assign memfont[4023] = 1'd0;
    assign memfont[4024] = 1'd0;
    assign memfont[4025] = 1'd0;
    assign memfont[4026] = 1'd0;
    assign memfont[4027] = 1'd0;
    assign memfont[4028] = 1'd0;
    assign memfont[4029] = 1'd1;
    assign memfont[4030] = 1'd1;
    assign memfont[4031] = 1'd0;
    assign memfont[4032] = 1'd0;
    assign memfont[4033] = 1'd1;
    assign memfont[4034] = 1'd1;
    assign memfont[4035] = 1'd0;
    assign memfont[4036] = 1'd0;
    assign memfont[4037] = 1'd0;
    assign memfont[4038] = 1'd1;
    assign memfont[4039] = 1'd1;
    assign memfont[4040] = 1'd0;
    assign memfont[4041] = 1'd0;
    assign memfont[4042] = 1'd0;
    assign memfont[4043] = 1'd0;
    assign memfont[4044] = 1'd0;
    assign memfont[4045] = 1'd0;
    assign memfont[4046] = 1'd0;
    assign memfont[4047] = 1'd0;
    assign memfont[4048] = 1'd0;
    assign memfont[4049] = 1'd0;
    assign memfont[4050] = 1'd0;
    assign memfont[4051] = 1'd0;
    assign memfont[4052] = 1'd1;
    assign memfont[4053] = 1'd1;
    assign memfont[4054] = 1'd1;
    assign memfont[4055] = 1'd0;
    assign memfont[4056] = 1'd0;
    assign memfont[4057] = 1'd0;
    assign memfont[4058] = 1'd0;
    assign memfont[4059] = 1'd0;
    assign memfont[4060] = 1'd0;
    assign memfont[4061] = 1'd1;
    assign memfont[4062] = 1'd1;
    assign memfont[4063] = 1'd0;
    assign memfont[4064] = 1'd0;
    assign memfont[4065] = 1'd0;
    assign memfont[4066] = 1'd0;
    assign memfont[4067] = 1'd0;
    assign memfont[4068] = 1'd0;
    assign memfont[4069] = 1'd1;
    assign memfont[4070] = 1'd1;
    assign memfont[4071] = 1'd0;
    assign memfont[4072] = 1'd0;
    assign memfont[4073] = 1'd0;
    assign memfont[4074] = 1'd0;
    assign memfont[4075] = 1'd0;
    assign memfont[4076] = 1'd0;
    assign memfont[4077] = 1'd1;
    assign memfont[4078] = 1'd1;
    assign memfont[4079] = 1'd0;
    assign memfont[4080] = 1'd0;
    assign memfont[4081] = 1'd0;
    assign memfont[4082] = 1'd0;
    assign memfont[4083] = 1'd1;
    assign memfont[4084] = 1'd1;
    assign memfont[4085] = 1'd0;
    assign memfont[4086] = 1'd0;
    assign memfont[4087] = 1'd1;
    assign memfont[4088] = 1'd1;
    assign memfont[4089] = 1'd0;
    assign memfont[4090] = 1'd0;
    assign memfont[4091] = 1'd0;
    assign memfont[4092] = 1'd0;
    assign memfont[4093] = 1'd1;
    assign memfont[4094] = 1'd1;
    assign memfont[4095] = 1'd1;
    assign memfont[4096] = 1'd1;
    assign memfont[4097] = 1'd0;
    assign memfont[4098] = 1'd0;
    assign memfont[4099] = 1'd1;
    assign memfont[4100] = 1'd1;
    assign memfont[4101] = 1'd1;
    assign memfont[4102] = 1'd0;
    assign memfont[4103] = 1'd0;
    assign memfont[4104] = 1'd0;
    assign memfont[4105] = 1'd0;
    assign memfont[4106] = 1'd0;
    assign memfont[4107] = 1'd0;
    assign memfont[4108] = 1'd1;
    assign memfont[4109] = 1'd1;
    assign memfont[4110] = 1'd1;
    assign memfont[4111] = 1'd1;
    assign memfont[4112] = 1'd0;
    assign memfont[4113] = 1'd0;
    assign memfont[4114] = 1'd0;
    assign memfont[4115] = 1'd0;
    assign memfont[4116] = 1'd0;
    assign memfont[4117] = 1'd0;
    assign memfont[4118] = 1'd0;
    assign memfont[4119] = 1'd0;
    assign memfont[4120] = 1'd0;
    assign memfont[4121] = 1'd1;
    assign memfont[4122] = 1'd1;
    assign memfont[4123] = 1'd0;
    assign memfont[4124] = 1'd0;
    assign memfont[4125] = 1'd0;
    assign memfont[4126] = 1'd0;
    assign memfont[4127] = 1'd0;
    assign memfont[4128] = 1'd0;
    assign memfont[4129] = 1'd0;
    assign memfont[4130] = 1'd0;
    assign memfont[4131] = 1'd1;
    assign memfont[4132] = 1'd1;
    assign memfont[4133] = 1'd1;
    assign memfont[4134] = 1'd0;
    assign memfont[4135] = 1'd0;
    assign memfont[4136] = 1'd0;
    assign memfont[4137] = 1'd0;
    assign memfont[4138] = 1'd0;
    assign memfont[4139] = 1'd0;
    assign memfont[4140] = 1'd0;
    assign memfont[4141] = 1'd0;
    assign memfont[4142] = 1'd0;
    assign memfont[4143] = 1'd0;
    assign memfont[4144] = 1'd0;
    assign memfont[4145] = 1'd1;
    assign memfont[4146] = 1'd1;
    assign memfont[4147] = 1'd0;
    assign memfont[4148] = 1'd0;
    assign memfont[4149] = 1'd0;
    assign memfont[4150] = 1'd0;
    assign memfont[4151] = 1'd0;
    assign memfont[4152] = 1'd0;
    assign memfont[4153] = 1'd1;
    assign memfont[4154] = 1'd1;
    assign memfont[4155] = 1'd0;
    assign memfont[4156] = 1'd0;
    assign memfont[4157] = 1'd0;
    assign memfont[4158] = 1'd0;
    assign memfont[4159] = 1'd0;
    assign memfont[4160] = 1'd0;
    assign memfont[4161] = 1'd1;
    assign memfont[4162] = 1'd1;
    assign memfont[4163] = 1'd0;
    assign memfont[4164] = 1'd0;
    assign memfont[4165] = 1'd1;
    assign memfont[4166] = 1'd1;
    assign memfont[4167] = 1'd1;
    assign memfont[4168] = 1'd1;
    assign memfont[4169] = 1'd1;
    assign memfont[4170] = 1'd1;
    assign memfont[4171] = 1'd1;
    assign memfont[4172] = 1'd1;
    assign memfont[4173] = 1'd1;
    assign memfont[4174] = 1'd1;
    assign memfont[4175] = 1'd0;
    assign memfont[4176] = 1'd0;
    assign memfont[4177] = 1'd0;
    assign memfont[4178] = 1'd1;
    assign memfont[4179] = 1'd1;
    assign memfont[4180] = 1'd1;
    assign memfont[4181] = 1'd1;
    assign memfont[4182] = 1'd1;
    assign memfont[4183] = 1'd1;
    assign memfont[4184] = 1'd1;
    assign memfont[4185] = 1'd1;
    assign memfont[4186] = 1'd0;
    assign memfont[4187] = 1'd0;
    assign memfont[4188] = 1'd0;
    assign memfont[4189] = 1'd1;
    assign memfont[4190] = 1'd1;
    assign memfont[4191] = 1'd0;
    assign memfont[4192] = 1'd0;
    assign memfont[4193] = 1'd0;
    assign memfont[4194] = 1'd0;
    assign memfont[4195] = 1'd0;
    assign memfont[4196] = 1'd0;
    assign memfont[4197] = 1'd1;
    assign memfont[4198] = 1'd1;
    assign memfont[4199] = 1'd0;
    assign memfont[4200] = 1'd0;
    assign memfont[4201] = 1'd1;
    assign memfont[4202] = 1'd1;
    assign memfont[4203] = 1'd0;
    assign memfont[4204] = 1'd0;
    assign memfont[4205] = 1'd0;
    assign memfont[4206] = 1'd0;
    assign memfont[4207] = 1'd0;
    assign memfont[4208] = 1'd0;
    assign memfont[4209] = 1'd1;
    assign memfont[4210] = 1'd1;
    assign memfont[4211] = 1'd0;
    assign memfont[4212] = 1'd0;
    assign memfont[4213] = 1'd1;
    assign memfont[4214] = 1'd1;
    assign memfont[4215] = 1'd0;
    assign memfont[4216] = 1'd0;
    assign memfont[4217] = 1'd0;
    assign memfont[4218] = 1'd0;
    assign memfont[4219] = 1'd0;
    assign memfont[4220] = 1'd1;
    assign memfont[4221] = 1'd1;
    assign memfont[4222] = 1'd1;
    assign memfont[4223] = 1'd0;
    assign memfont[4224] = 1'd0;
    assign memfont[4225] = 1'd1;
    assign memfont[4226] = 1'd1;
    assign memfont[4227] = 1'd0;
    assign memfont[4228] = 1'd0;
    assign memfont[4229] = 1'd0;
    assign memfont[4230] = 1'd0;
    assign memfont[4231] = 1'd0;
    assign memfont[4232] = 1'd0;
    assign memfont[4233] = 1'd0;
    assign memfont[4234] = 1'd0;
    assign memfont[4235] = 1'd0;
    assign memfont[4236] = 1'd0;
    assign memfont[4237] = 1'd1;
    assign memfont[4238] = 1'd1;
    assign memfont[4239] = 1'd0;
    assign memfont[4240] = 1'd0;
    assign memfont[4241] = 1'd0;
    assign memfont[4242] = 1'd0;
    assign memfont[4243] = 1'd0;
    assign memfont[4244] = 1'd0;
    assign memfont[4245] = 1'd0;
    assign memfont[4246] = 1'd0;
    assign memfont[4247] = 1'd0;
    assign memfont[4248] = 1'd0;
    assign memfont[4249] = 1'd1;
    assign memfont[4250] = 1'd1;
    assign memfont[4251] = 1'd0;
    assign memfont[4252] = 1'd0;
    assign memfont[4253] = 1'd0;
    assign memfont[4254] = 1'd0;
    assign memfont[4255] = 1'd0;
    assign memfont[4256] = 1'd0;
    assign memfont[4257] = 1'd1;
    assign memfont[4258] = 1'd1;
    assign memfont[4259] = 1'd0;
    assign memfont[4260] = 1'd0;
    assign memfont[4261] = 1'd1;
    assign memfont[4262] = 1'd1;
    assign memfont[4263] = 1'd0;
    assign memfont[4264] = 1'd0;
    assign memfont[4265] = 1'd0;
    assign memfont[4266] = 1'd0;
    assign memfont[4267] = 1'd0;
    assign memfont[4268] = 1'd0;
    assign memfont[4269] = 1'd1;
    assign memfont[4270] = 1'd1;
    assign memfont[4271] = 1'd0;
    assign memfont[4272] = 1'd0;
    assign memfont[4273] = 1'd0;
    assign memfont[4274] = 1'd0;
    assign memfont[4275] = 1'd0;
    assign memfont[4276] = 1'd0;
    assign memfont[4277] = 1'd1;
    assign memfont[4278] = 1'd1;
    assign memfont[4279] = 1'd0;
    assign memfont[4280] = 1'd0;
    assign memfont[4281] = 1'd0;
    assign memfont[4282] = 1'd0;
    assign memfont[4283] = 1'd0;
    assign memfont[4284] = 1'd0;
    assign memfont[4285] = 1'd1;
    assign memfont[4286] = 1'd1;
    assign memfont[4287] = 1'd0;
    assign memfont[4288] = 1'd0;
    assign memfont[4289] = 1'd0;
    assign memfont[4290] = 1'd0;
    assign memfont[4291] = 1'd0;
    assign memfont[4292] = 1'd1;
    assign memfont[4293] = 1'd1;
    assign memfont[4294] = 1'd0;
    assign memfont[4295] = 1'd0;
    assign memfont[4296] = 1'd0;
    assign memfont[4297] = 1'd1;
    assign memfont[4298] = 1'd1;
    assign memfont[4299] = 1'd0;
    assign memfont[4300] = 1'd0;
    assign memfont[4301] = 1'd0;
    assign memfont[4302] = 1'd1;
    assign memfont[4303] = 1'd1;
    assign memfont[4304] = 1'd1;
    assign memfont[4305] = 1'd0;
    assign memfont[4306] = 1'd0;
    assign memfont[4307] = 1'd0;
    assign memfont[4308] = 1'd0;
    assign memfont[4309] = 1'd1;
    assign memfont[4310] = 1'd1;
    assign memfont[4311] = 1'd0;
    assign memfont[4312] = 1'd0;
    assign memfont[4313] = 1'd0;
    assign memfont[4314] = 1'd0;
    assign memfont[4315] = 1'd0;
    assign memfont[4316] = 1'd0;
    assign memfont[4317] = 1'd0;
    assign memfont[4318] = 1'd0;
    assign memfont[4319] = 1'd0;
    assign memfont[4320] = 1'd0;
    assign memfont[4321] = 1'd1;
    assign memfont[4322] = 1'd1;
    assign memfont[4323] = 1'd0;
    assign memfont[4324] = 1'd1;
    assign memfont[4325] = 1'd1;
    assign memfont[4326] = 1'd1;
    assign memfont[4327] = 1'd1;
    assign memfont[4328] = 1'd0;
    assign memfont[4329] = 1'd1;
    assign memfont[4330] = 1'd1;
    assign memfont[4331] = 1'd0;
    assign memfont[4332] = 1'd0;
    assign memfont[4333] = 1'd1;
    assign memfont[4334] = 1'd1;
    assign memfont[4335] = 1'd0;
    assign memfont[4336] = 1'd0;
    assign memfont[4337] = 1'd0;
    assign memfont[4338] = 1'd1;
    assign memfont[4339] = 1'd1;
    assign memfont[4340] = 1'd0;
    assign memfont[4341] = 1'd1;
    assign memfont[4342] = 1'd1;
    assign memfont[4343] = 1'd0;
    assign memfont[4344] = 1'd0;
    assign memfont[4345] = 1'd1;
    assign memfont[4346] = 1'd1;
    assign memfont[4347] = 1'd0;
    assign memfont[4348] = 1'd0;
    assign memfont[4349] = 1'd0;
    assign memfont[4350] = 1'd0;
    assign memfont[4351] = 1'd0;
    assign memfont[4352] = 1'd0;
    assign memfont[4353] = 1'd1;
    assign memfont[4354] = 1'd1;
    assign memfont[4355] = 1'd0;
    assign memfont[4356] = 1'd0;
    assign memfont[4357] = 1'd1;
    assign memfont[4358] = 1'd1;
    assign memfont[4359] = 1'd0;
    assign memfont[4360] = 1'd0;
    assign memfont[4361] = 1'd0;
    assign memfont[4362] = 1'd0;
    assign memfont[4363] = 1'd0;
    assign memfont[4364] = 1'd0;
    assign memfont[4365] = 1'd0;
    assign memfont[4366] = 1'd0;
    assign memfont[4367] = 1'd0;
    assign memfont[4368] = 1'd0;
    assign memfont[4369] = 1'd1;
    assign memfont[4370] = 1'd1;
    assign memfont[4371] = 1'd0;
    assign memfont[4372] = 1'd0;
    assign memfont[4373] = 1'd0;
    assign memfont[4374] = 1'd1;
    assign memfont[4375] = 1'd1;
    assign memfont[4376] = 1'd0;
    assign memfont[4377] = 1'd1;
    assign memfont[4378] = 1'd1;
    assign memfont[4379] = 1'd0;
    assign memfont[4380] = 1'd0;
    assign memfont[4381] = 1'd1;
    assign memfont[4382] = 1'd1;
    assign memfont[4383] = 1'd0;
    assign memfont[4384] = 1'd0;
    assign memfont[4385] = 1'd0;
    assign memfont[4386] = 1'd0;
    assign memfont[4387] = 1'd1;
    assign memfont[4388] = 1'd1;
    assign memfont[4389] = 1'd0;
    assign memfont[4390] = 1'd0;
    assign memfont[4391] = 1'd0;
    assign memfont[4392] = 1'd0;
    assign memfont[4393] = 1'd1;
    assign memfont[4394] = 1'd1;
    assign memfont[4395] = 1'd0;
    assign memfont[4396] = 1'd0;
    assign memfont[4397] = 1'd0;
    assign memfont[4398] = 1'd0;
    assign memfont[4399] = 1'd0;
    assign memfont[4400] = 1'd0;
    assign memfont[4401] = 1'd1;
    assign memfont[4402] = 1'd1;
    assign memfont[4403] = 1'd0;
    assign memfont[4404] = 1'd0;
    assign memfont[4405] = 1'd0;
    assign memfont[4406] = 1'd0;
    assign memfont[4407] = 1'd0;
    assign memfont[4408] = 1'd0;
    assign memfont[4409] = 1'd1;
    assign memfont[4410] = 1'd1;
    assign memfont[4411] = 1'd0;
    assign memfont[4412] = 1'd0;
    assign memfont[4413] = 1'd0;
    assign memfont[4414] = 1'd0;
    assign memfont[4415] = 1'd0;
    assign memfont[4416] = 1'd0;
    assign memfont[4417] = 1'd1;
    assign memfont[4418] = 1'd1;
    assign memfont[4419] = 1'd0;
    assign memfont[4420] = 1'd0;
    assign memfont[4421] = 1'd0;
    assign memfont[4422] = 1'd0;
    assign memfont[4423] = 1'd0;
    assign memfont[4424] = 1'd0;
    assign memfont[4425] = 1'd1;
    assign memfont[4426] = 1'd1;
    assign memfont[4427] = 1'd0;
    assign memfont[4428] = 1'd0;
    assign memfont[4429] = 1'd0;
    assign memfont[4430] = 1'd0;
    assign memfont[4431] = 1'd1;
    assign memfont[4432] = 1'd1;
    assign memfont[4433] = 1'd0;
    assign memfont[4434] = 1'd1;
    assign memfont[4435] = 1'd1;
    assign memfont[4436] = 1'd0;
    assign memfont[4437] = 1'd0;
    assign memfont[4438] = 1'd0;
    assign memfont[4439] = 1'd0;
    assign memfont[4440] = 1'd0;
    assign memfont[4441] = 1'd1;
    assign memfont[4442] = 1'd1;
    assign memfont[4443] = 1'd1;
    assign memfont[4444] = 1'd1;
    assign memfont[4445] = 1'd0;
    assign memfont[4446] = 1'd0;
    assign memfont[4447] = 1'd1;
    assign memfont[4448] = 1'd1;
    assign memfont[4449] = 1'd1;
    assign memfont[4450] = 1'd0;
    assign memfont[4451] = 1'd0;
    assign memfont[4452] = 1'd0;
    assign memfont[4453] = 1'd0;
    assign memfont[4454] = 1'd0;
    assign memfont[4455] = 1'd1;
    assign memfont[4456] = 1'd1;
    assign memfont[4457] = 1'd0;
    assign memfont[4458] = 1'd0;
    assign memfont[4459] = 1'd1;
    assign memfont[4460] = 1'd1;
    assign memfont[4461] = 1'd0;
    assign memfont[4462] = 1'd0;
    assign memfont[4463] = 1'd0;
    assign memfont[4464] = 1'd0;
    assign memfont[4465] = 1'd0;
    assign memfont[4466] = 1'd0;
    assign memfont[4467] = 1'd0;
    assign memfont[4468] = 1'd0;
    assign memfont[4469] = 1'd1;
    assign memfont[4470] = 1'd1;
    assign memfont[4471] = 1'd0;
    assign memfont[4472] = 1'd0;
    assign memfont[4473] = 1'd0;
    assign memfont[4474] = 1'd0;
    assign memfont[4475] = 1'd0;
    assign memfont[4476] = 1'd0;
    assign memfont[4477] = 1'd0;
    assign memfont[4478] = 1'd0;
    assign memfont[4479] = 1'd1;
    assign memfont[4480] = 1'd1;
    assign memfont[4481] = 1'd0;
    assign memfont[4482] = 1'd0;
    assign memfont[4483] = 1'd0;
    assign memfont[4484] = 1'd0;
    assign memfont[4485] = 1'd0;
    assign memfont[4486] = 1'd0;
    assign memfont[4487] = 1'd0;
    assign memfont[4488] = 1'd0;
    assign memfont[4489] = 1'd0;
    assign memfont[4490] = 1'd0;
    assign memfont[4491] = 1'd0;
    assign memfont[4492] = 1'd0;
    assign memfont[4493] = 1'd1;
    assign memfont[4494] = 1'd0;
    assign memfont[4495] = 1'd0;
    assign memfont[4496] = 1'd0;
    assign memfont[4497] = 1'd0;
    assign memfont[4498] = 1'd0;
    assign memfont[4499] = 1'd0;
    assign memfont[4500] = 1'd0;
    assign memfont[4501] = 1'd1;
    assign memfont[4502] = 1'd1;
    assign memfont[4503] = 1'd1;
    assign memfont[4504] = 1'd0;
    assign memfont[4505] = 1'd0;
    assign memfont[4506] = 1'd0;
    assign memfont[4507] = 1'd0;
    assign memfont[4508] = 1'd1;
    assign memfont[4509] = 1'd1;
    assign memfont[4510] = 1'd1;
    assign memfont[4511] = 1'd0;
    assign memfont[4512] = 1'd0;
    assign memfont[4513] = 1'd1;
    assign memfont[4514] = 1'd1;
    assign memfont[4515] = 1'd1;
    assign memfont[4516] = 1'd1;
    assign memfont[4517] = 1'd1;
    assign memfont[4518] = 1'd1;
    assign memfont[4519] = 1'd1;
    assign memfont[4520] = 1'd1;
    assign memfont[4521] = 1'd1;
    assign memfont[4522] = 1'd1;
    assign memfont[4523] = 1'd0;
    assign memfont[4524] = 1'd0;
    assign memfont[4525] = 1'd1;
    assign memfont[4526] = 1'd1;
    assign memfont[4527] = 1'd1;
    assign memfont[4528] = 1'd0;
    assign memfont[4529] = 1'd0;
    assign memfont[4530] = 1'd0;
    assign memfont[4531] = 1'd0;
    assign memfont[4532] = 1'd1;
    assign memfont[4533] = 1'd1;
    assign memfont[4534] = 1'd0;
    assign memfont[4535] = 1'd0;
    assign memfont[4536] = 1'd0;
    assign memfont[4537] = 1'd1;
    assign memfont[4538] = 1'd1;
    assign memfont[4539] = 1'd0;
    assign memfont[4540] = 1'd0;
    assign memfont[4541] = 1'd0;
    assign memfont[4542] = 1'd0;
    assign memfont[4543] = 1'd0;
    assign memfont[4544] = 1'd0;
    assign memfont[4545] = 1'd1;
    assign memfont[4546] = 1'd1;
    assign memfont[4547] = 1'd0;
    assign memfont[4548] = 1'd0;
    assign memfont[4549] = 1'd1;
    assign memfont[4550] = 1'd1;
    assign memfont[4551] = 1'd1;
    assign memfont[4552] = 1'd0;
    assign memfont[4553] = 1'd0;
    assign memfont[4554] = 1'd0;
    assign memfont[4555] = 1'd0;
    assign memfont[4556] = 1'd0;
    assign memfont[4557] = 1'd1;
    assign memfont[4558] = 1'd1;
    assign memfont[4559] = 1'd0;
    assign memfont[4560] = 1'd0;
    assign memfont[4561] = 1'd1;
    assign memfont[4562] = 1'd1;
    assign memfont[4563] = 1'd0;
    assign memfont[4564] = 1'd0;
    assign memfont[4565] = 1'd0;
    assign memfont[4566] = 1'd0;
    assign memfont[4567] = 1'd0;
    assign memfont[4568] = 1'd1;
    assign memfont[4569] = 1'd1;
    assign memfont[4570] = 1'd0;
    assign memfont[4571] = 1'd0;
    assign memfont[4572] = 1'd0;
    assign memfont[4573] = 1'd1;
    assign memfont[4574] = 1'd1;
    assign memfont[4575] = 1'd0;
    assign memfont[4576] = 1'd0;
    assign memfont[4577] = 1'd0;
    assign memfont[4578] = 1'd0;
    assign memfont[4579] = 1'd0;
    assign memfont[4580] = 1'd0;
    assign memfont[4581] = 1'd0;
    assign memfont[4582] = 1'd0;
    assign memfont[4583] = 1'd0;
    assign memfont[4584] = 1'd0;
    assign memfont[4585] = 1'd1;
    assign memfont[4586] = 1'd1;
    assign memfont[4587] = 1'd0;
    assign memfont[4588] = 1'd0;
    assign memfont[4589] = 1'd0;
    assign memfont[4590] = 1'd0;
    assign memfont[4591] = 1'd0;
    assign memfont[4592] = 1'd0;
    assign memfont[4593] = 1'd0;
    assign memfont[4594] = 1'd0;
    assign memfont[4595] = 1'd0;
    assign memfont[4596] = 1'd0;
    assign memfont[4597] = 1'd1;
    assign memfont[4598] = 1'd1;
    assign memfont[4599] = 1'd1;
    assign memfont[4600] = 1'd0;
    assign memfont[4601] = 1'd0;
    assign memfont[4602] = 1'd0;
    assign memfont[4603] = 1'd0;
    assign memfont[4604] = 1'd0;
    assign memfont[4605] = 1'd1;
    assign memfont[4606] = 1'd1;
    assign memfont[4607] = 1'd0;
    assign memfont[4608] = 1'd0;
    assign memfont[4609] = 1'd1;
    assign memfont[4610] = 1'd1;
    assign memfont[4611] = 1'd0;
    assign memfont[4612] = 1'd0;
    assign memfont[4613] = 1'd0;
    assign memfont[4614] = 1'd0;
    assign memfont[4615] = 1'd0;
    assign memfont[4616] = 1'd0;
    assign memfont[4617] = 1'd1;
    assign memfont[4618] = 1'd1;
    assign memfont[4619] = 1'd0;
    assign memfont[4620] = 1'd0;
    assign memfont[4621] = 1'd0;
    assign memfont[4622] = 1'd0;
    assign memfont[4623] = 1'd0;
    assign memfont[4624] = 1'd0;
    assign memfont[4625] = 1'd1;
    assign memfont[4626] = 1'd1;
    assign memfont[4627] = 1'd0;
    assign memfont[4628] = 1'd0;
    assign memfont[4629] = 1'd0;
    assign memfont[4630] = 1'd0;
    assign memfont[4631] = 1'd0;
    assign memfont[4632] = 1'd0;
    assign memfont[4633] = 1'd1;
    assign memfont[4634] = 1'd1;
    assign memfont[4635] = 1'd0;
    assign memfont[4636] = 1'd0;
    assign memfont[4637] = 1'd0;
    assign memfont[4638] = 1'd0;
    assign memfont[4639] = 1'd0;
    assign memfont[4640] = 1'd1;
    assign memfont[4641] = 1'd1;
    assign memfont[4642] = 1'd0;
    assign memfont[4643] = 1'd0;
    assign memfont[4644] = 1'd0;
    assign memfont[4645] = 1'd1;
    assign memfont[4646] = 1'd1;
    assign memfont[4647] = 1'd0;
    assign memfont[4648] = 1'd0;
    assign memfont[4649] = 1'd0;
    assign memfont[4650] = 1'd0;
    assign memfont[4651] = 1'd1;
    assign memfont[4652] = 1'd1;
    assign memfont[4653] = 1'd0;
    assign memfont[4654] = 1'd0;
    assign memfont[4655] = 1'd0;
    assign memfont[4656] = 1'd0;
    assign memfont[4657] = 1'd1;
    assign memfont[4658] = 1'd1;
    assign memfont[4659] = 1'd0;
    assign memfont[4660] = 1'd0;
    assign memfont[4661] = 1'd0;
    assign memfont[4662] = 1'd0;
    assign memfont[4663] = 1'd0;
    assign memfont[4664] = 1'd0;
    assign memfont[4665] = 1'd0;
    assign memfont[4666] = 1'd0;
    assign memfont[4667] = 1'd0;
    assign memfont[4668] = 1'd0;
    assign memfont[4669] = 1'd1;
    assign memfont[4670] = 1'd1;
    assign memfont[4671] = 1'd0;
    assign memfont[4672] = 1'd1;
    assign memfont[4673] = 1'd1;
    assign memfont[4674] = 1'd1;
    assign memfont[4675] = 1'd0;
    assign memfont[4676] = 1'd0;
    assign memfont[4677] = 1'd1;
    assign memfont[4678] = 1'd1;
    assign memfont[4679] = 1'd0;
    assign memfont[4680] = 1'd0;
    assign memfont[4681] = 1'd1;
    assign memfont[4682] = 1'd1;
    assign memfont[4683] = 1'd0;
    assign memfont[4684] = 1'd0;
    assign memfont[4685] = 1'd0;
    assign memfont[4686] = 1'd0;
    assign memfont[4687] = 1'd1;
    assign memfont[4688] = 1'd1;
    assign memfont[4689] = 1'd1;
    assign memfont[4690] = 1'd1;
    assign memfont[4691] = 1'd0;
    assign memfont[4692] = 1'd0;
    assign memfont[4693] = 1'd1;
    assign memfont[4694] = 1'd1;
    assign memfont[4695] = 1'd0;
    assign memfont[4696] = 1'd0;
    assign memfont[4697] = 1'd0;
    assign memfont[4698] = 1'd0;
    assign memfont[4699] = 1'd0;
    assign memfont[4700] = 1'd1;
    assign memfont[4701] = 1'd1;
    assign memfont[4702] = 1'd1;
    assign memfont[4703] = 1'd0;
    assign memfont[4704] = 1'd0;
    assign memfont[4705] = 1'd1;
    assign memfont[4706] = 1'd1;
    assign memfont[4707] = 1'd0;
    assign memfont[4708] = 1'd0;
    assign memfont[4709] = 1'd0;
    assign memfont[4710] = 1'd0;
    assign memfont[4711] = 1'd0;
    assign memfont[4712] = 1'd0;
    assign memfont[4713] = 1'd0;
    assign memfont[4714] = 1'd0;
    assign memfont[4715] = 1'd0;
    assign memfont[4716] = 1'd0;
    assign memfont[4717] = 1'd1;
    assign memfont[4718] = 1'd1;
    assign memfont[4719] = 1'd0;
    assign memfont[4720] = 1'd0;
    assign memfont[4721] = 1'd0;
    assign memfont[4722] = 1'd1;
    assign memfont[4723] = 1'd1;
    assign memfont[4724] = 1'd1;
    assign memfont[4725] = 1'd1;
    assign memfont[4726] = 1'd1;
    assign memfont[4727] = 1'd0;
    assign memfont[4728] = 1'd0;
    assign memfont[4729] = 1'd1;
    assign memfont[4730] = 1'd1;
    assign memfont[4731] = 1'd0;
    assign memfont[4732] = 1'd0;
    assign memfont[4733] = 1'd0;
    assign memfont[4734] = 1'd0;
    assign memfont[4735] = 1'd1;
    assign memfont[4736] = 1'd1;
    assign memfont[4737] = 1'd0;
    assign memfont[4738] = 1'd0;
    assign memfont[4739] = 1'd0;
    assign memfont[4740] = 1'd0;
    assign memfont[4741] = 1'd1;
    assign memfont[4742] = 1'd1;
    assign memfont[4743] = 1'd0;
    assign memfont[4744] = 1'd0;
    assign memfont[4745] = 1'd0;
    assign memfont[4746] = 1'd0;
    assign memfont[4747] = 1'd0;
    assign memfont[4748] = 1'd0;
    assign memfont[4749] = 1'd1;
    assign memfont[4750] = 1'd1;
    assign memfont[4751] = 1'd0;
    assign memfont[4752] = 1'd0;
    assign memfont[4753] = 1'd0;
    assign memfont[4754] = 1'd0;
    assign memfont[4755] = 1'd0;
    assign memfont[4756] = 1'd0;
    assign memfont[4757] = 1'd1;
    assign memfont[4758] = 1'd1;
    assign memfont[4759] = 1'd0;
    assign memfont[4760] = 1'd0;
    assign memfont[4761] = 1'd0;
    assign memfont[4762] = 1'd0;
    assign memfont[4763] = 1'd0;
    assign memfont[4764] = 1'd0;
    assign memfont[4765] = 1'd1;
    assign memfont[4766] = 1'd1;
    assign memfont[4767] = 1'd0;
    assign memfont[4768] = 1'd0;
    assign memfont[4769] = 1'd0;
    assign memfont[4770] = 1'd0;
    assign memfont[4771] = 1'd0;
    assign memfont[4772] = 1'd0;
    assign memfont[4773] = 1'd1;
    assign memfont[4774] = 1'd1;
    assign memfont[4775] = 1'd0;
    assign memfont[4776] = 1'd0;
    assign memfont[4777] = 1'd0;
    assign memfont[4778] = 1'd0;
    assign memfont[4779] = 1'd0;
    assign memfont[4780] = 1'd1;
    assign memfont[4781] = 1'd1;
    assign memfont[4782] = 1'd1;
    assign memfont[4783] = 1'd1;
    assign memfont[4784] = 1'd0;
    assign memfont[4785] = 1'd0;
    assign memfont[4786] = 1'd0;
    assign memfont[4787] = 1'd0;
    assign memfont[4788] = 1'd0;
    assign memfont[4789] = 1'd0;
    assign memfont[4790] = 1'd1;
    assign memfont[4791] = 1'd1;
    assign memfont[4792] = 1'd1;
    assign memfont[4793] = 1'd0;
    assign memfont[4794] = 1'd0;
    assign memfont[4795] = 1'd1;
    assign memfont[4796] = 1'd1;
    assign memfont[4797] = 1'd1;
    assign memfont[4798] = 1'd0;
    assign memfont[4799] = 1'd0;
    assign memfont[4800] = 1'd0;
    assign memfont[4801] = 1'd0;
    assign memfont[4802] = 1'd1;
    assign memfont[4803] = 1'd1;
    assign memfont[4804] = 1'd1;
    assign memfont[4805] = 1'd0;
    assign memfont[4806] = 1'd0;
    assign memfont[4807] = 1'd1;
    assign memfont[4808] = 1'd1;
    assign memfont[4809] = 1'd0;
    assign memfont[4810] = 1'd0;
    assign memfont[4811] = 1'd0;
    assign memfont[4812] = 1'd0;
    assign memfont[4813] = 1'd0;
    assign memfont[4814] = 1'd0;
    assign memfont[4815] = 1'd0;
    assign memfont[4816] = 1'd0;
    assign memfont[4817] = 1'd1;
    assign memfont[4818] = 1'd1;
    assign memfont[4819] = 1'd0;
    assign memfont[4820] = 1'd0;
    assign memfont[4821] = 1'd0;
    assign memfont[4822] = 1'd0;
    assign memfont[4823] = 1'd0;
    assign memfont[4824] = 1'd0;
    assign memfont[4825] = 1'd0;
    assign memfont[4826] = 1'd1;
    assign memfont[4827] = 1'd1;
    assign memfont[4828] = 1'd0;
    assign memfont[4829] = 1'd0;
    assign memfont[4830] = 1'd0;
    assign memfont[4831] = 1'd0;
    assign memfont[4832] = 1'd0;
    assign memfont[4833] = 1'd0;
    assign memfont[4834] = 1'd0;
    assign memfont[4835] = 1'd0;
    assign memfont[4836] = 1'd0;
    assign memfont[4837] = 1'd0;
    assign memfont[4838] = 1'd0;
    assign memfont[4839] = 1'd0;
    assign memfont[4840] = 1'd0;
    assign memfont[4841] = 1'd0;
    assign memfont[4842] = 1'd0;
    assign memfont[4843] = 1'd0;
    assign memfont[4844] = 1'd0;
    assign memfont[4845] = 1'd0;
    assign memfont[4846] = 1'd0;
    assign memfont[4847] = 1'd0;
    assign memfont[4848] = 1'd0;
    assign memfont[4849] = 1'd1;
    assign memfont[4850] = 1'd1;
    assign memfont[4851] = 1'd1;
    assign memfont[4852] = 1'd1;
    assign memfont[4853] = 1'd1;
    assign memfont[4854] = 1'd1;
    assign memfont[4855] = 1'd1;
    assign memfont[4856] = 1'd1;
    assign memfont[4857] = 1'd1;
    assign memfont[4858] = 1'd1;
    assign memfont[4859] = 1'd0;
    assign memfont[4860] = 1'd0;
    assign memfont[4861] = 1'd1;
    assign memfont[4862] = 1'd1;
    assign memfont[4863] = 1'd1;
    assign memfont[4864] = 1'd1;
    assign memfont[4865] = 1'd1;
    assign memfont[4866] = 1'd1;
    assign memfont[4867] = 1'd1;
    assign memfont[4868] = 1'd1;
    assign memfont[4869] = 1'd1;
    assign memfont[4870] = 1'd1;
    assign memfont[4871] = 1'd0;
    assign memfont[4872] = 1'd0;
    assign memfont[4873] = 1'd1;
    assign memfont[4874] = 1'd1;
    assign memfont[4875] = 1'd0;
    assign memfont[4876] = 1'd0;
    assign memfont[4877] = 1'd0;
    assign memfont[4878] = 1'd0;
    assign memfont[4879] = 1'd0;
    assign memfont[4880] = 1'd1;
    assign memfont[4881] = 1'd1;
    assign memfont[4882] = 1'd1;
    assign memfont[4883] = 1'd0;
    assign memfont[4884] = 1'd0;
    assign memfont[4885] = 1'd1;
    assign memfont[4886] = 1'd1;
    assign memfont[4887] = 1'd0;
    assign memfont[4888] = 1'd0;
    assign memfont[4889] = 1'd0;
    assign memfont[4890] = 1'd0;
    assign memfont[4891] = 1'd0;
    assign memfont[4892] = 1'd1;
    assign memfont[4893] = 1'd1;
    assign memfont[4894] = 1'd1;
    assign memfont[4895] = 1'd0;
    assign memfont[4896] = 1'd0;
    assign memfont[4897] = 1'd0;
    assign memfont[4898] = 1'd1;
    assign memfont[4899] = 1'd1;
    assign memfont[4900] = 1'd0;
    assign memfont[4901] = 1'd0;
    assign memfont[4902] = 1'd0;
    assign memfont[4903] = 1'd0;
    assign memfont[4904] = 1'd1;
    assign memfont[4905] = 1'd1;
    assign memfont[4906] = 1'd1;
    assign memfont[4907] = 1'd0;
    assign memfont[4908] = 1'd0;
    assign memfont[4909] = 1'd1;
    assign memfont[4910] = 1'd1;
    assign memfont[4911] = 1'd0;
    assign memfont[4912] = 1'd0;
    assign memfont[4913] = 1'd0;
    assign memfont[4914] = 1'd0;
    assign memfont[4915] = 1'd1;
    assign memfont[4916] = 1'd1;
    assign memfont[4917] = 1'd1;
    assign memfont[4918] = 1'd0;
    assign memfont[4919] = 1'd0;
    assign memfont[4920] = 1'd0;
    assign memfont[4921] = 1'd1;
    assign memfont[4922] = 1'd1;
    assign memfont[4923] = 1'd0;
    assign memfont[4924] = 1'd0;
    assign memfont[4925] = 1'd0;
    assign memfont[4926] = 1'd0;
    assign memfont[4927] = 1'd0;
    assign memfont[4928] = 1'd0;
    assign memfont[4929] = 1'd0;
    assign memfont[4930] = 1'd0;
    assign memfont[4931] = 1'd0;
    assign memfont[4932] = 1'd0;
    assign memfont[4933] = 1'd1;
    assign memfont[4934] = 1'd1;
    assign memfont[4935] = 1'd0;
    assign memfont[4936] = 1'd0;
    assign memfont[4937] = 1'd0;
    assign memfont[4938] = 1'd0;
    assign memfont[4939] = 1'd0;
    assign memfont[4940] = 1'd0;
    assign memfont[4941] = 1'd0;
    assign memfont[4942] = 1'd0;
    assign memfont[4943] = 1'd0;
    assign memfont[4944] = 1'd0;
    assign memfont[4945] = 1'd0;
    assign memfont[4946] = 1'd1;
    assign memfont[4947] = 1'd1;
    assign memfont[4948] = 1'd0;
    assign memfont[4949] = 1'd0;
    assign memfont[4950] = 1'd0;
    assign memfont[4951] = 1'd0;
    assign memfont[4952] = 1'd1;
    assign memfont[4953] = 1'd1;
    assign memfont[4954] = 1'd1;
    assign memfont[4955] = 1'd0;
    assign memfont[4956] = 1'd0;
    assign memfont[4957] = 1'd1;
    assign memfont[4958] = 1'd1;
    assign memfont[4959] = 1'd0;
    assign memfont[4960] = 1'd0;
    assign memfont[4961] = 1'd0;
    assign memfont[4962] = 1'd0;
    assign memfont[4963] = 1'd0;
    assign memfont[4964] = 1'd0;
    assign memfont[4965] = 1'd1;
    assign memfont[4966] = 1'd1;
    assign memfont[4967] = 1'd0;
    assign memfont[4968] = 1'd0;
    assign memfont[4969] = 1'd0;
    assign memfont[4970] = 1'd0;
    assign memfont[4971] = 1'd0;
    assign memfont[4972] = 1'd0;
    assign memfont[4973] = 1'd1;
    assign memfont[4974] = 1'd1;
    assign memfont[4975] = 1'd0;
    assign memfont[4976] = 1'd0;
    assign memfont[4977] = 1'd0;
    assign memfont[4978] = 1'd0;
    assign memfont[4979] = 1'd0;
    assign memfont[4980] = 1'd0;
    assign memfont[4981] = 1'd1;
    assign memfont[4982] = 1'd1;
    assign memfont[4983] = 1'd1;
    assign memfont[4984] = 1'd0;
    assign memfont[4985] = 1'd0;
    assign memfont[4986] = 1'd0;
    assign memfont[4987] = 1'd0;
    assign memfont[4988] = 1'd1;
    assign memfont[4989] = 1'd1;
    assign memfont[4990] = 1'd0;
    assign memfont[4991] = 1'd0;
    assign memfont[4992] = 1'd0;
    assign memfont[4993] = 1'd1;
    assign memfont[4994] = 1'd1;
    assign memfont[4995] = 1'd0;
    assign memfont[4996] = 1'd0;
    assign memfont[4997] = 1'd0;
    assign memfont[4998] = 1'd0;
    assign memfont[4999] = 1'd1;
    assign memfont[5000] = 1'd1;
    assign memfont[5001] = 1'd1;
    assign memfont[5002] = 1'd0;
    assign memfont[5003] = 1'd0;
    assign memfont[5004] = 1'd0;
    assign memfont[5005] = 1'd1;
    assign memfont[5006] = 1'd1;
    assign memfont[5007] = 1'd0;
    assign memfont[5008] = 1'd0;
    assign memfont[5009] = 1'd0;
    assign memfont[5010] = 1'd0;
    assign memfont[5011] = 1'd0;
    assign memfont[5012] = 1'd0;
    assign memfont[5013] = 1'd0;
    assign memfont[5014] = 1'd0;
    assign memfont[5015] = 1'd0;
    assign memfont[5016] = 1'd0;
    assign memfont[5017] = 1'd1;
    assign memfont[5018] = 1'd1;
    assign memfont[5019] = 1'd0;
    assign memfont[5020] = 1'd0;
    assign memfont[5021] = 1'd1;
    assign memfont[5022] = 1'd1;
    assign memfont[5023] = 1'd0;
    assign memfont[5024] = 1'd0;
    assign memfont[5025] = 1'd1;
    assign memfont[5026] = 1'd1;
    assign memfont[5027] = 1'd0;
    assign memfont[5028] = 1'd0;
    assign memfont[5029] = 1'd1;
    assign memfont[5030] = 1'd1;
    assign memfont[5031] = 1'd0;
    assign memfont[5032] = 1'd0;
    assign memfont[5033] = 1'd0;
    assign memfont[5034] = 1'd0;
    assign memfont[5035] = 1'd1;
    assign memfont[5036] = 1'd1;
    assign memfont[5037] = 1'd1;
    assign memfont[5038] = 1'd1;
    assign memfont[5039] = 1'd0;
    assign memfont[5040] = 1'd0;
    assign memfont[5041] = 1'd1;
    assign memfont[5042] = 1'd1;
    assign memfont[5043] = 1'd1;
    assign memfont[5044] = 1'd0;
    assign memfont[5045] = 1'd0;
    assign memfont[5046] = 1'd0;
    assign memfont[5047] = 1'd0;
    assign memfont[5048] = 1'd1;
    assign memfont[5049] = 1'd1;
    assign memfont[5050] = 1'd0;
    assign memfont[5051] = 1'd0;
    assign memfont[5052] = 1'd0;
    assign memfont[5053] = 1'd1;
    assign memfont[5054] = 1'd1;
    assign memfont[5055] = 1'd0;
    assign memfont[5056] = 1'd0;
    assign memfont[5057] = 1'd0;
    assign memfont[5058] = 1'd0;
    assign memfont[5059] = 1'd0;
    assign memfont[5060] = 1'd0;
    assign memfont[5061] = 1'd0;
    assign memfont[5062] = 1'd0;
    assign memfont[5063] = 1'd0;
    assign memfont[5064] = 1'd0;
    assign memfont[5065] = 1'd1;
    assign memfont[5066] = 1'd1;
    assign memfont[5067] = 1'd1;
    assign memfont[5068] = 1'd0;
    assign memfont[5069] = 1'd0;
    assign memfont[5070] = 1'd0;
    assign memfont[5071] = 1'd1;
    assign memfont[5072] = 1'd1;
    assign memfont[5073] = 1'd1;
    assign memfont[5074] = 1'd0;
    assign memfont[5075] = 1'd0;
    assign memfont[5076] = 1'd0;
    assign memfont[5077] = 1'd1;
    assign memfont[5078] = 1'd1;
    assign memfont[5079] = 1'd0;
    assign memfont[5080] = 1'd0;
    assign memfont[5081] = 1'd0;
    assign memfont[5082] = 1'd0;
    assign memfont[5083] = 1'd0;
    assign memfont[5084] = 1'd1;
    assign memfont[5085] = 1'd1;
    assign memfont[5086] = 1'd0;
    assign memfont[5087] = 1'd0;
    assign memfont[5088] = 1'd0;
    assign memfont[5089] = 1'd1;
    assign memfont[5090] = 1'd1;
    assign memfont[5091] = 1'd0;
    assign memfont[5092] = 1'd0;
    assign memfont[5093] = 1'd0;
    assign memfont[5094] = 1'd0;
    assign memfont[5095] = 1'd0;
    assign memfont[5096] = 1'd1;
    assign memfont[5097] = 1'd1;
    assign memfont[5098] = 1'd1;
    assign memfont[5099] = 1'd0;
    assign memfont[5100] = 1'd0;
    assign memfont[5101] = 1'd0;
    assign memfont[5102] = 1'd0;
    assign memfont[5103] = 1'd0;
    assign memfont[5104] = 1'd0;
    assign memfont[5105] = 1'd1;
    assign memfont[5106] = 1'd1;
    assign memfont[5107] = 1'd0;
    assign memfont[5108] = 1'd0;
    assign memfont[5109] = 1'd0;
    assign memfont[5110] = 1'd0;
    assign memfont[5111] = 1'd0;
    assign memfont[5112] = 1'd0;
    assign memfont[5113] = 1'd1;
    assign memfont[5114] = 1'd1;
    assign memfont[5115] = 1'd0;
    assign memfont[5116] = 1'd0;
    assign memfont[5117] = 1'd0;
    assign memfont[5118] = 1'd0;
    assign memfont[5119] = 1'd0;
    assign memfont[5120] = 1'd1;
    assign memfont[5121] = 1'd1;
    assign memfont[5122] = 1'd1;
    assign memfont[5123] = 1'd0;
    assign memfont[5124] = 1'd0;
    assign memfont[5125] = 1'd0;
    assign memfont[5126] = 1'd0;
    assign memfont[5127] = 1'd0;
    assign memfont[5128] = 1'd1;
    assign memfont[5129] = 1'd1;
    assign memfont[5130] = 1'd1;
    assign memfont[5131] = 1'd1;
    assign memfont[5132] = 1'd0;
    assign memfont[5133] = 1'd0;
    assign memfont[5134] = 1'd0;
    assign memfont[5135] = 1'd0;
    assign memfont[5136] = 1'd0;
    assign memfont[5137] = 1'd0;
    assign memfont[5138] = 1'd1;
    assign memfont[5139] = 1'd1;
    assign memfont[5140] = 1'd0;
    assign memfont[5141] = 1'd0;
    assign memfont[5142] = 1'd0;
    assign memfont[5143] = 1'd1;
    assign memfont[5144] = 1'd1;
    assign memfont[5145] = 1'd1;
    assign memfont[5146] = 1'd0;
    assign memfont[5147] = 1'd0;
    assign memfont[5148] = 1'd0;
    assign memfont[5149] = 1'd0;
    assign memfont[5150] = 1'd1;
    assign memfont[5151] = 1'd1;
    assign memfont[5152] = 1'd0;
    assign memfont[5153] = 1'd0;
    assign memfont[5154] = 1'd0;
    assign memfont[5155] = 1'd0;
    assign memfont[5156] = 1'd1;
    assign memfont[5157] = 1'd1;
    assign memfont[5158] = 1'd0;
    assign memfont[5159] = 1'd0;
    assign memfont[5160] = 1'd0;
    assign memfont[5161] = 1'd0;
    assign memfont[5162] = 1'd0;
    assign memfont[5163] = 1'd0;
    assign memfont[5164] = 1'd0;
    assign memfont[5165] = 1'd1;
    assign memfont[5166] = 1'd1;
    assign memfont[5167] = 1'd0;
    assign memfont[5168] = 1'd0;
    assign memfont[5169] = 1'd0;
    assign memfont[5170] = 1'd0;
    assign memfont[5171] = 1'd0;
    assign memfont[5172] = 1'd0;
    assign memfont[5173] = 1'd0;
    assign memfont[5174] = 1'd1;
    assign memfont[5175] = 1'd1;
    assign memfont[5176] = 1'd0;
    assign memfont[5177] = 1'd0;
    assign memfont[5178] = 1'd0;
    assign memfont[5179] = 1'd0;
    assign memfont[5180] = 1'd0;
    assign memfont[5181] = 1'd0;
    assign memfont[5182] = 1'd0;
    assign memfont[5183] = 1'd0;
    assign memfont[5184] = 1'd0;
    assign memfont[5185] = 1'd0;
    assign memfont[5186] = 1'd0;
    assign memfont[5187] = 1'd0;
    assign memfont[5188] = 1'd0;
    assign memfont[5189] = 1'd0;
    assign memfont[5190] = 1'd0;
    assign memfont[5191] = 1'd0;
    assign memfont[5192] = 1'd0;
    assign memfont[5193] = 1'd0;
    assign memfont[5194] = 1'd0;
    assign memfont[5195] = 1'd0;
    assign memfont[5196] = 1'd0;
    assign memfont[5197] = 1'd0;
    assign memfont[5198] = 1'd0;
    assign memfont[5199] = 1'd0;
    assign memfont[5200] = 1'd0;
    assign memfont[5201] = 1'd0;
    assign memfont[5202] = 1'd0;
    assign memfont[5203] = 1'd0;
    assign memfont[5204] = 1'd0;
    assign memfont[5205] = 1'd0;
    assign memfont[5206] = 1'd0;
    assign memfont[5207] = 1'd0;
    assign memfont[5208] = 1'd0;
    assign memfont[5209] = 1'd0;
    assign memfont[5210] = 1'd0;
    assign memfont[5211] = 1'd0;
    assign memfont[5212] = 1'd0;
    assign memfont[5213] = 1'd0;
    assign memfont[5214] = 1'd0;
    assign memfont[5215] = 1'd0;
    assign memfont[5216] = 1'd0;
    assign memfont[5217] = 1'd0;
    assign memfont[5218] = 1'd0;
    assign memfont[5219] = 1'd0;
    assign memfont[5220] = 1'd0;
    assign memfont[5221] = 1'd1;
    assign memfont[5222] = 1'd1;
    assign memfont[5223] = 1'd0;
    assign memfont[5224] = 1'd0;
    assign memfont[5225] = 1'd0;
    assign memfont[5226] = 1'd0;
    assign memfont[5227] = 1'd0;
    assign memfont[5228] = 1'd0;
    assign memfont[5229] = 1'd1;
    assign memfont[5230] = 1'd1;
    assign memfont[5231] = 1'd0;
    assign memfont[5232] = 1'd0;
    assign memfont[5233] = 1'd1;
    assign memfont[5234] = 1'd1;
    assign memfont[5235] = 1'd0;
    assign memfont[5236] = 1'd0;
    assign memfont[5237] = 1'd0;
    assign memfont[5238] = 1'd0;
    assign memfont[5239] = 1'd1;
    assign memfont[5240] = 1'd1;
    assign memfont[5241] = 1'd1;
    assign memfont[5242] = 1'd0;
    assign memfont[5243] = 1'd0;
    assign memfont[5244] = 1'd0;
    assign memfont[5245] = 1'd0;
    assign memfont[5246] = 1'd1;
    assign memfont[5247] = 1'd1;
    assign memfont[5248] = 1'd1;
    assign memfont[5249] = 1'd0;
    assign memfont[5250] = 1'd0;
    assign memfont[5251] = 1'd0;
    assign memfont[5252] = 1'd1;
    assign memfont[5253] = 1'd1;
    assign memfont[5254] = 1'd0;
    assign memfont[5255] = 1'd0;
    assign memfont[5256] = 1'd0;
    assign memfont[5257] = 1'd1;
    assign memfont[5258] = 1'd1;
    assign memfont[5259] = 1'd0;
    assign memfont[5260] = 1'd0;
    assign memfont[5261] = 1'd0;
    assign memfont[5262] = 1'd1;
    assign memfont[5263] = 1'd1;
    assign memfont[5264] = 1'd1;
    assign memfont[5265] = 1'd0;
    assign memfont[5266] = 1'd0;
    assign memfont[5267] = 1'd0;
    assign memfont[5268] = 1'd0;
    assign memfont[5269] = 1'd1;
    assign memfont[5270] = 1'd1;
    assign memfont[5271] = 1'd0;
    assign memfont[5272] = 1'd0;
    assign memfont[5273] = 1'd0;
    assign memfont[5274] = 1'd0;
    assign memfont[5275] = 1'd0;
    assign memfont[5276] = 1'd0;
    assign memfont[5277] = 1'd0;
    assign memfont[5278] = 1'd0;
    assign memfont[5279] = 1'd0;
    assign memfont[5280] = 1'd0;
    assign memfont[5281] = 1'd1;
    assign memfont[5282] = 1'd1;
    assign memfont[5283] = 1'd0;
    assign memfont[5284] = 1'd0;
    assign memfont[5285] = 1'd0;
    assign memfont[5286] = 1'd0;
    assign memfont[5287] = 1'd0;
    assign memfont[5288] = 1'd0;
    assign memfont[5289] = 1'd0;
    assign memfont[5290] = 1'd0;
    assign memfont[5291] = 1'd0;
    assign memfont[5292] = 1'd0;
    assign memfont[5293] = 1'd0;
    assign memfont[5294] = 1'd1;
    assign memfont[5295] = 1'd1;
    assign memfont[5296] = 1'd1;
    assign memfont[5297] = 1'd0;
    assign memfont[5298] = 1'd0;
    assign memfont[5299] = 1'd0;
    assign memfont[5300] = 1'd1;
    assign memfont[5301] = 1'd1;
    assign memfont[5302] = 1'd1;
    assign memfont[5303] = 1'd0;
    assign memfont[5304] = 1'd0;
    assign memfont[5305] = 1'd1;
    assign memfont[5306] = 1'd1;
    assign memfont[5307] = 1'd0;
    assign memfont[5308] = 1'd0;
    assign memfont[5309] = 1'd0;
    assign memfont[5310] = 1'd0;
    assign memfont[5311] = 1'd0;
    assign memfont[5312] = 1'd0;
    assign memfont[5313] = 1'd1;
    assign memfont[5314] = 1'd1;
    assign memfont[5315] = 1'd0;
    assign memfont[5316] = 1'd0;
    assign memfont[5317] = 1'd0;
    assign memfont[5318] = 1'd0;
    assign memfont[5319] = 1'd0;
    assign memfont[5320] = 1'd0;
    assign memfont[5321] = 1'd1;
    assign memfont[5322] = 1'd1;
    assign memfont[5323] = 1'd0;
    assign memfont[5324] = 1'd0;
    assign memfont[5325] = 1'd0;
    assign memfont[5326] = 1'd0;
    assign memfont[5327] = 1'd0;
    assign memfont[5328] = 1'd0;
    assign memfont[5329] = 1'd0;
    assign memfont[5330] = 1'd1;
    assign memfont[5331] = 1'd1;
    assign memfont[5332] = 1'd1;
    assign memfont[5333] = 1'd0;
    assign memfont[5334] = 1'd0;
    assign memfont[5335] = 1'd1;
    assign memfont[5336] = 1'd1;
    assign memfont[5337] = 1'd1;
    assign memfont[5338] = 1'd0;
    assign memfont[5339] = 1'd0;
    assign memfont[5340] = 1'd0;
    assign memfont[5341] = 1'd1;
    assign memfont[5342] = 1'd1;
    assign memfont[5343] = 1'd0;
    assign memfont[5344] = 1'd0;
    assign memfont[5345] = 1'd0;
    assign memfont[5346] = 1'd0;
    assign memfont[5347] = 1'd0;
    assign memfont[5348] = 1'd1;
    assign memfont[5349] = 1'd1;
    assign memfont[5350] = 1'd0;
    assign memfont[5351] = 1'd0;
    assign memfont[5352] = 1'd0;
    assign memfont[5353] = 1'd1;
    assign memfont[5354] = 1'd1;
    assign memfont[5355] = 1'd0;
    assign memfont[5356] = 1'd0;
    assign memfont[5357] = 1'd0;
    assign memfont[5358] = 1'd0;
    assign memfont[5359] = 1'd0;
    assign memfont[5360] = 1'd0;
    assign memfont[5361] = 1'd0;
    assign memfont[5362] = 1'd0;
    assign memfont[5363] = 1'd0;
    assign memfont[5364] = 1'd0;
    assign memfont[5365] = 1'd1;
    assign memfont[5366] = 1'd1;
    assign memfont[5367] = 1'd0;
    assign memfont[5368] = 1'd0;
    assign memfont[5369] = 1'd1;
    assign memfont[5370] = 1'd1;
    assign memfont[5371] = 1'd0;
    assign memfont[5372] = 1'd0;
    assign memfont[5373] = 1'd1;
    assign memfont[5374] = 1'd1;
    assign memfont[5375] = 1'd0;
    assign memfont[5376] = 1'd0;
    assign memfont[5377] = 1'd1;
    assign memfont[5378] = 1'd1;
    assign memfont[5379] = 1'd0;
    assign memfont[5380] = 1'd0;
    assign memfont[5381] = 1'd0;
    assign memfont[5382] = 1'd0;
    assign memfont[5383] = 1'd1;
    assign memfont[5384] = 1'd1;
    assign memfont[5385] = 1'd1;
    assign memfont[5386] = 1'd1;
    assign memfont[5387] = 1'd0;
    assign memfont[5388] = 1'd0;
    assign memfont[5389] = 1'd0;
    assign memfont[5390] = 1'd1;
    assign memfont[5391] = 1'd1;
    assign memfont[5392] = 1'd1;
    assign memfont[5393] = 1'd0;
    assign memfont[5394] = 1'd0;
    assign memfont[5395] = 1'd1;
    assign memfont[5396] = 1'd1;
    assign memfont[5397] = 1'd1;
    assign memfont[5398] = 1'd0;
    assign memfont[5399] = 1'd0;
    assign memfont[5400] = 1'd0;
    assign memfont[5401] = 1'd1;
    assign memfont[5402] = 1'd1;
    assign memfont[5403] = 1'd0;
    assign memfont[5404] = 1'd0;
    assign memfont[5405] = 1'd0;
    assign memfont[5406] = 1'd0;
    assign memfont[5407] = 1'd0;
    assign memfont[5408] = 1'd0;
    assign memfont[5409] = 1'd0;
    assign memfont[5410] = 1'd0;
    assign memfont[5411] = 1'd0;
    assign memfont[5412] = 1'd0;
    assign memfont[5413] = 1'd0;
    assign memfont[5414] = 1'd1;
    assign memfont[5415] = 1'd1;
    assign memfont[5416] = 1'd1;
    assign memfont[5417] = 1'd0;
    assign memfont[5418] = 1'd0;
    assign memfont[5419] = 1'd1;
    assign memfont[5420] = 1'd1;
    assign memfont[5421] = 1'd1;
    assign memfont[5422] = 1'd0;
    assign memfont[5423] = 1'd0;
    assign memfont[5424] = 1'd0;
    assign memfont[5425] = 1'd1;
    assign memfont[5426] = 1'd1;
    assign memfont[5427] = 1'd0;
    assign memfont[5428] = 1'd0;
    assign memfont[5429] = 1'd0;
    assign memfont[5430] = 1'd0;
    assign memfont[5431] = 1'd0;
    assign memfont[5432] = 1'd1;
    assign memfont[5433] = 1'd1;
    assign memfont[5434] = 1'd0;
    assign memfont[5435] = 1'd0;
    assign memfont[5436] = 1'd0;
    assign memfont[5437] = 1'd1;
    assign memfont[5438] = 1'd1;
    assign memfont[5439] = 1'd1;
    assign memfont[5440] = 1'd0;
    assign memfont[5441] = 1'd0;
    assign memfont[5442] = 1'd0;
    assign memfont[5443] = 1'd0;
    assign memfont[5444] = 1'd1;
    assign memfont[5445] = 1'd1;
    assign memfont[5446] = 1'd0;
    assign memfont[5447] = 1'd0;
    assign memfont[5448] = 1'd0;
    assign memfont[5449] = 1'd0;
    assign memfont[5450] = 1'd0;
    assign memfont[5451] = 1'd0;
    assign memfont[5452] = 1'd0;
    assign memfont[5453] = 1'd1;
    assign memfont[5454] = 1'd1;
    assign memfont[5455] = 1'd0;
    assign memfont[5456] = 1'd0;
    assign memfont[5457] = 1'd0;
    assign memfont[5458] = 1'd0;
    assign memfont[5459] = 1'd0;
    assign memfont[5460] = 1'd0;
    assign memfont[5461] = 1'd0;
    assign memfont[5462] = 1'd1;
    assign memfont[5463] = 1'd1;
    assign memfont[5464] = 1'd0;
    assign memfont[5465] = 1'd0;
    assign memfont[5466] = 1'd0;
    assign memfont[5467] = 1'd1;
    assign memfont[5468] = 1'd1;
    assign memfont[5469] = 1'd1;
    assign memfont[5470] = 1'd0;
    assign memfont[5471] = 1'd0;
    assign memfont[5472] = 1'd0;
    assign memfont[5473] = 1'd0;
    assign memfont[5474] = 1'd0;
    assign memfont[5475] = 1'd0;
    assign memfont[5476] = 1'd1;
    assign memfont[5477] = 1'd1;
    assign memfont[5478] = 1'd1;
    assign memfont[5479] = 1'd0;
    assign memfont[5480] = 1'd0;
    assign memfont[5481] = 1'd0;
    assign memfont[5482] = 1'd0;
    assign memfont[5483] = 1'd0;
    assign memfont[5484] = 1'd0;
    assign memfont[5485] = 1'd0;
    assign memfont[5486] = 1'd1;
    assign memfont[5487] = 1'd1;
    assign memfont[5488] = 1'd0;
    assign memfont[5489] = 1'd0;
    assign memfont[5490] = 1'd0;
    assign memfont[5491] = 1'd1;
    assign memfont[5492] = 1'd1;
    assign memfont[5493] = 1'd1;
    assign memfont[5494] = 1'd0;
    assign memfont[5495] = 1'd0;
    assign memfont[5496] = 1'd0;
    assign memfont[5497] = 1'd1;
    assign memfont[5498] = 1'd1;
    assign memfont[5499] = 1'd1;
    assign memfont[5500] = 1'd0;
    assign memfont[5501] = 1'd0;
    assign memfont[5502] = 1'd0;
    assign memfont[5503] = 1'd0;
    assign memfont[5504] = 1'd1;
    assign memfont[5505] = 1'd1;
    assign memfont[5506] = 1'd0;
    assign memfont[5507] = 1'd0;
    assign memfont[5508] = 1'd0;
    assign memfont[5509] = 1'd0;
    assign memfont[5510] = 1'd0;
    assign memfont[5511] = 1'd0;
    assign memfont[5512] = 1'd0;
    assign memfont[5513] = 1'd1;
    assign memfont[5514] = 1'd1;
    assign memfont[5515] = 1'd0;
    assign memfont[5516] = 1'd0;
    assign memfont[5517] = 1'd0;
    assign memfont[5518] = 1'd0;
    assign memfont[5519] = 1'd0;
    assign memfont[5520] = 1'd0;
    assign memfont[5521] = 1'd1;
    assign memfont[5522] = 1'd1;
    assign memfont[5523] = 1'd0;
    assign memfont[5524] = 1'd0;
    assign memfont[5525] = 1'd0;
    assign memfont[5526] = 1'd0;
    assign memfont[5527] = 1'd0;
    assign memfont[5528] = 1'd0;
    assign memfont[5529] = 1'd0;
    assign memfont[5530] = 1'd0;
    assign memfont[5531] = 1'd0;
    assign memfont[5532] = 1'd0;
    assign memfont[5533] = 1'd0;
    assign memfont[5534] = 1'd0;
    assign memfont[5535] = 1'd0;
    assign memfont[5536] = 1'd1;
    assign memfont[5537] = 1'd1;
    assign memfont[5538] = 1'd1;
    assign memfont[5539] = 1'd0;
    assign memfont[5540] = 1'd0;
    assign memfont[5541] = 1'd0;
    assign memfont[5542] = 1'd0;
    assign memfont[5543] = 1'd0;
    assign memfont[5544] = 1'd0;
    assign memfont[5545] = 1'd0;
    assign memfont[5546] = 1'd0;
    assign memfont[5547] = 1'd0;
    assign memfont[5548] = 1'd0;
    assign memfont[5549] = 1'd0;
    assign memfont[5550] = 1'd0;
    assign memfont[5551] = 1'd0;
    assign memfont[5552] = 1'd0;
    assign memfont[5553] = 1'd0;
    assign memfont[5554] = 1'd0;
    assign memfont[5555] = 1'd0;
    assign memfont[5556] = 1'd0;
    assign memfont[5557] = 1'd0;
    assign memfont[5558] = 1'd0;
    assign memfont[5559] = 1'd0;
    assign memfont[5560] = 1'd0;
    assign memfont[5561] = 1'd0;
    assign memfont[5562] = 1'd0;
    assign memfont[5563] = 1'd0;
    assign memfont[5564] = 1'd0;
    assign memfont[5565] = 1'd0;
    assign memfont[5566] = 1'd0;
    assign memfont[5567] = 1'd0;
    assign memfont[5568] = 1'd0;
    assign memfont[5569] = 1'd1;
    assign memfont[5570] = 1'd1;
    assign memfont[5571] = 1'd0;
    assign memfont[5572] = 1'd0;
    assign memfont[5573] = 1'd0;
    assign memfont[5574] = 1'd0;
    assign memfont[5575] = 1'd0;
    assign memfont[5576] = 1'd0;
    assign memfont[5577] = 1'd1;
    assign memfont[5578] = 1'd1;
    assign memfont[5579] = 1'd0;
    assign memfont[5580] = 1'd0;
    assign memfont[5581] = 1'd1;
    assign memfont[5582] = 1'd1;
    assign memfont[5583] = 1'd1;
    assign memfont[5584] = 1'd1;
    assign memfont[5585] = 1'd1;
    assign memfont[5586] = 1'd1;
    assign memfont[5587] = 1'd1;
    assign memfont[5588] = 1'd1;
    assign memfont[5589] = 1'd1;
    assign memfont[5590] = 1'd0;
    assign memfont[5591] = 1'd0;
    assign memfont[5592] = 1'd0;
    assign memfont[5593] = 1'd0;
    assign memfont[5594] = 1'd0;
    assign memfont[5595] = 1'd1;
    assign memfont[5596] = 1'd1;
    assign memfont[5597] = 1'd1;
    assign memfont[5598] = 1'd1;
    assign memfont[5599] = 1'd1;
    assign memfont[5600] = 1'd1;
    assign memfont[5601] = 1'd0;
    assign memfont[5602] = 1'd0;
    assign memfont[5603] = 1'd0;
    assign memfont[5604] = 1'd0;
    assign memfont[5605] = 1'd1;
    assign memfont[5606] = 1'd1;
    assign memfont[5607] = 1'd1;
    assign memfont[5608] = 1'd1;
    assign memfont[5609] = 1'd1;
    assign memfont[5610] = 1'd1;
    assign memfont[5611] = 1'd1;
    assign memfont[5612] = 1'd0;
    assign memfont[5613] = 1'd0;
    assign memfont[5614] = 1'd0;
    assign memfont[5615] = 1'd0;
    assign memfont[5616] = 1'd0;
    assign memfont[5617] = 1'd1;
    assign memfont[5618] = 1'd1;
    assign memfont[5619] = 1'd1;
    assign memfont[5620] = 1'd1;
    assign memfont[5621] = 1'd1;
    assign memfont[5622] = 1'd1;
    assign memfont[5623] = 1'd1;
    assign memfont[5624] = 1'd1;
    assign memfont[5625] = 1'd1;
    assign memfont[5626] = 1'd1;
    assign memfont[5627] = 1'd0;
    assign memfont[5628] = 1'd0;
    assign memfont[5629] = 1'd1;
    assign memfont[5630] = 1'd1;
    assign memfont[5631] = 1'd0;
    assign memfont[5632] = 1'd0;
    assign memfont[5633] = 1'd0;
    assign memfont[5634] = 1'd0;
    assign memfont[5635] = 1'd0;
    assign memfont[5636] = 1'd0;
    assign memfont[5637] = 1'd0;
    assign memfont[5638] = 1'd0;
    assign memfont[5639] = 1'd0;
    assign memfont[5640] = 1'd0;
    assign memfont[5641] = 1'd0;
    assign memfont[5642] = 1'd0;
    assign memfont[5643] = 1'd1;
    assign memfont[5644] = 1'd1;
    assign memfont[5645] = 1'd1;
    assign memfont[5646] = 1'd1;
    assign memfont[5647] = 1'd1;
    assign memfont[5648] = 1'd1;
    assign memfont[5649] = 1'd1;
    assign memfont[5650] = 1'd1;
    assign memfont[5651] = 1'd0;
    assign memfont[5652] = 1'd0;
    assign memfont[5653] = 1'd1;
    assign memfont[5654] = 1'd1;
    assign memfont[5655] = 1'd0;
    assign memfont[5656] = 1'd0;
    assign memfont[5657] = 1'd0;
    assign memfont[5658] = 1'd0;
    assign memfont[5659] = 1'd0;
    assign memfont[5660] = 1'd0;
    assign memfont[5661] = 1'd1;
    assign memfont[5662] = 1'd1;
    assign memfont[5663] = 1'd0;
    assign memfont[5664] = 1'd0;
    assign memfont[5665] = 1'd0;
    assign memfont[5666] = 1'd0;
    assign memfont[5667] = 1'd0;
    assign memfont[5668] = 1'd0;
    assign memfont[5669] = 1'd1;
    assign memfont[5670] = 1'd1;
    assign memfont[5671] = 1'd0;
    assign memfont[5672] = 1'd0;
    assign memfont[5673] = 1'd0;
    assign memfont[5674] = 1'd0;
    assign memfont[5675] = 1'd0;
    assign memfont[5676] = 1'd0;
    assign memfont[5677] = 1'd0;
    assign memfont[5678] = 1'd0;
    assign memfont[5679] = 1'd1;
    assign memfont[5680] = 1'd1;
    assign memfont[5681] = 1'd1;
    assign memfont[5682] = 1'd1;
    assign memfont[5683] = 1'd1;
    assign memfont[5684] = 1'd1;
    assign memfont[5685] = 1'd0;
    assign memfont[5686] = 1'd0;
    assign memfont[5687] = 1'd0;
    assign memfont[5688] = 1'd0;
    assign memfont[5689] = 1'd1;
    assign memfont[5690] = 1'd1;
    assign memfont[5691] = 1'd0;
    assign memfont[5692] = 1'd0;
    assign memfont[5693] = 1'd0;
    assign memfont[5694] = 1'd0;
    assign memfont[5695] = 1'd0;
    assign memfont[5696] = 1'd1;
    assign memfont[5697] = 1'd1;
    assign memfont[5698] = 1'd1;
    assign memfont[5699] = 1'd0;
    assign memfont[5700] = 1'd0;
    assign memfont[5701] = 1'd1;
    assign memfont[5702] = 1'd1;
    assign memfont[5703] = 1'd1;
    assign memfont[5704] = 1'd1;
    assign memfont[5705] = 1'd1;
    assign memfont[5706] = 1'd1;
    assign memfont[5707] = 1'd1;
    assign memfont[5708] = 1'd1;
    assign memfont[5709] = 1'd1;
    assign memfont[5710] = 1'd1;
    assign memfont[5711] = 1'd0;
    assign memfont[5712] = 1'd0;
    assign memfont[5713] = 1'd1;
    assign memfont[5714] = 1'd1;
    assign memfont[5715] = 1'd0;
    assign memfont[5716] = 1'd0;
    assign memfont[5717] = 1'd1;
    assign memfont[5718] = 1'd1;
    assign memfont[5719] = 1'd0;
    assign memfont[5720] = 1'd0;
    assign memfont[5721] = 1'd1;
    assign memfont[5722] = 1'd1;
    assign memfont[5723] = 1'd0;
    assign memfont[5724] = 1'd0;
    assign memfont[5725] = 1'd1;
    assign memfont[5726] = 1'd1;
    assign memfont[5727] = 1'd0;
    assign memfont[5728] = 1'd0;
    assign memfont[5729] = 1'd0;
    assign memfont[5730] = 1'd0;
    assign memfont[5731] = 1'd0;
    assign memfont[5732] = 1'd1;
    assign memfont[5733] = 1'd1;
    assign memfont[5734] = 1'd1;
    assign memfont[5735] = 1'd0;
    assign memfont[5736] = 1'd0;
    assign memfont[5737] = 1'd0;
    assign memfont[5738] = 1'd0;
    assign memfont[5739] = 1'd1;
    assign memfont[5740] = 1'd1;
    assign memfont[5741] = 1'd1;
    assign memfont[5742] = 1'd1;
    assign memfont[5743] = 1'd1;
    assign memfont[5744] = 1'd1;
    assign memfont[5745] = 1'd0;
    assign memfont[5746] = 1'd0;
    assign memfont[5747] = 1'd0;
    assign memfont[5748] = 1'd0;
    assign memfont[5749] = 1'd1;
    assign memfont[5750] = 1'd1;
    assign memfont[5751] = 1'd0;
    assign memfont[5752] = 1'd0;
    assign memfont[5753] = 1'd0;
    assign memfont[5754] = 1'd0;
    assign memfont[5755] = 1'd0;
    assign memfont[5756] = 1'd0;
    assign memfont[5757] = 1'd0;
    assign memfont[5758] = 1'd0;
    assign memfont[5759] = 1'd0;
    assign memfont[5760] = 1'd0;
    assign memfont[5761] = 1'd0;
    assign memfont[5762] = 1'd0;
    assign memfont[5763] = 1'd1;
    assign memfont[5764] = 1'd1;
    assign memfont[5765] = 1'd1;
    assign memfont[5766] = 1'd1;
    assign memfont[5767] = 1'd1;
    assign memfont[5768] = 1'd1;
    assign memfont[5769] = 1'd1;
    assign memfont[5770] = 1'd0;
    assign memfont[5771] = 1'd0;
    assign memfont[5772] = 1'd0;
    assign memfont[5773] = 1'd1;
    assign memfont[5774] = 1'd1;
    assign memfont[5775] = 1'd0;
    assign memfont[5776] = 1'd0;
    assign memfont[5777] = 1'd0;
    assign memfont[5778] = 1'd0;
    assign memfont[5779] = 1'd0;
    assign memfont[5780] = 1'd1;
    assign memfont[5781] = 1'd1;
    assign memfont[5782] = 1'd1;
    assign memfont[5783] = 1'd0;
    assign memfont[5784] = 1'd0;
    assign memfont[5785] = 1'd0;
    assign memfont[5786] = 1'd1;
    assign memfont[5787] = 1'd1;
    assign memfont[5788] = 1'd1;
    assign memfont[5789] = 1'd1;
    assign memfont[5790] = 1'd1;
    assign memfont[5791] = 1'd1;
    assign memfont[5792] = 1'd1;
    assign memfont[5793] = 1'd0;
    assign memfont[5794] = 1'd0;
    assign memfont[5795] = 1'd0;
    assign memfont[5796] = 1'd0;
    assign memfont[5797] = 1'd0;
    assign memfont[5798] = 1'd0;
    assign memfont[5799] = 1'd0;
    assign memfont[5800] = 1'd0;
    assign memfont[5801] = 1'd1;
    assign memfont[5802] = 1'd1;
    assign memfont[5803] = 1'd0;
    assign memfont[5804] = 1'd0;
    assign memfont[5805] = 1'd0;
    assign memfont[5806] = 1'd0;
    assign memfont[5807] = 1'd0;
    assign memfont[5808] = 1'd0;
    assign memfont[5809] = 1'd0;
    assign memfont[5810] = 1'd1;
    assign memfont[5811] = 1'd1;
    assign memfont[5812] = 1'd1;
    assign memfont[5813] = 1'd1;
    assign memfont[5814] = 1'd1;
    assign memfont[5815] = 1'd1;
    assign memfont[5816] = 1'd1;
    assign memfont[5817] = 1'd1;
    assign memfont[5818] = 1'd0;
    assign memfont[5819] = 1'd0;
    assign memfont[5820] = 1'd0;
    assign memfont[5821] = 1'd0;
    assign memfont[5822] = 1'd0;
    assign memfont[5823] = 1'd0;
    assign memfont[5824] = 1'd0;
    assign memfont[5825] = 1'd1;
    assign memfont[5826] = 1'd1;
    assign memfont[5827] = 1'd0;
    assign memfont[5828] = 1'd0;
    assign memfont[5829] = 1'd0;
    assign memfont[5830] = 1'd0;
    assign memfont[5831] = 1'd0;
    assign memfont[5832] = 1'd0;
    assign memfont[5833] = 1'd0;
    assign memfont[5834] = 1'd1;
    assign memfont[5835] = 1'd1;
    assign memfont[5836] = 1'd0;
    assign memfont[5837] = 1'd0;
    assign memfont[5838] = 1'd0;
    assign memfont[5839] = 1'd1;
    assign memfont[5840] = 1'd1;
    assign memfont[5841] = 1'd1;
    assign memfont[5842] = 1'd0;
    assign memfont[5843] = 1'd0;
    assign memfont[5844] = 1'd0;
    assign memfont[5845] = 1'd1;
    assign memfont[5846] = 1'd1;
    assign memfont[5847] = 1'd0;
    assign memfont[5848] = 1'd0;
    assign memfont[5849] = 1'd0;
    assign memfont[5850] = 1'd0;
    assign memfont[5851] = 1'd0;
    assign memfont[5852] = 1'd1;
    assign memfont[5853] = 1'd1;
    assign memfont[5854] = 1'd1;
    assign memfont[5855] = 1'd0;
    assign memfont[5856] = 1'd0;
    assign memfont[5857] = 1'd0;
    assign memfont[5858] = 1'd0;
    assign memfont[5859] = 1'd0;
    assign memfont[5860] = 1'd0;
    assign memfont[5861] = 1'd1;
    assign memfont[5862] = 1'd1;
    assign memfont[5863] = 1'd0;
    assign memfont[5864] = 1'd0;
    assign memfont[5865] = 1'd0;
    assign memfont[5866] = 1'd0;
    assign memfont[5867] = 1'd0;
    assign memfont[5868] = 1'd0;
    assign memfont[5869] = 1'd1;
    assign memfont[5870] = 1'd1;
    assign memfont[5871] = 1'd1;
    assign memfont[5872] = 1'd1;
    assign memfont[5873] = 1'd1;
    assign memfont[5874] = 1'd1;
    assign memfont[5875] = 1'd1;
    assign memfont[5876] = 1'd1;
    assign memfont[5877] = 1'd1;
    assign memfont[5878] = 1'd1;
    assign memfont[5879] = 1'd0;
    assign memfont[5880] = 1'd0;
    assign memfont[5881] = 1'd0;
    assign memfont[5882] = 1'd0;
    assign memfont[5883] = 1'd0;
    assign memfont[5884] = 1'd1;
    assign memfont[5885] = 1'd1;
    assign memfont[5886] = 1'd1;
    assign memfont[5887] = 1'd0;
    assign memfont[5888] = 1'd0;
    assign memfont[5889] = 1'd0;
    assign memfont[5890] = 1'd0;
    assign memfont[5891] = 1'd0;
    assign memfont[5892] = 1'd0;
    assign memfont[5893] = 1'd0;
    assign memfont[5894] = 1'd0;
    assign memfont[5895] = 1'd0;
    assign memfont[5896] = 1'd0;
    assign memfont[5897] = 1'd0;
    assign memfont[5898] = 1'd0;
    assign memfont[5899] = 1'd0;
    assign memfont[5900] = 1'd0;
    assign memfont[5901] = 1'd0;
    assign memfont[5902] = 1'd0;
    assign memfont[5903] = 1'd0;
    assign memfont[5904] = 1'd0;
    assign memfont[5905] = 1'd0;
    assign memfont[5906] = 1'd0;
    assign memfont[5907] = 1'd0;
    assign memfont[5908] = 1'd0;
    assign memfont[5909] = 1'd0;
    assign memfont[5910] = 1'd0;
    assign memfont[5911] = 1'd0;
    assign memfont[5912] = 1'd0;
    assign memfont[5913] = 1'd0;
    assign memfont[5914] = 1'd0;
    assign memfont[5915] = 1'd0;
    assign memfont[5916] = 1'd1;
    assign memfont[5917] = 1'd1;
    assign memfont[5918] = 1'd1;
    assign memfont[5919] = 1'd0;
    assign memfont[5920] = 1'd0;
    assign memfont[5921] = 1'd0;
    assign memfont[5922] = 1'd0;
    assign memfont[5923] = 1'd0;
    assign memfont[5924] = 1'd0;
    assign memfont[5925] = 1'd1;
    assign memfont[5926] = 1'd1;
    assign memfont[5927] = 1'd1;
    assign memfont[5928] = 1'd0;
    assign memfont[5929] = 1'd1;
    assign memfont[5930] = 1'd1;
    assign memfont[5931] = 1'd1;
    assign memfont[5932] = 1'd1;
    assign memfont[5933] = 1'd1;
    assign memfont[5934] = 1'd1;
    assign memfont[5935] = 1'd0;
    assign memfont[5936] = 1'd0;
    assign memfont[5937] = 1'd0;
    assign memfont[5938] = 1'd0;
    assign memfont[5939] = 1'd0;
    assign memfont[5940] = 1'd0;
    assign memfont[5941] = 1'd0;
    assign memfont[5942] = 1'd0;
    assign memfont[5943] = 1'd0;
    assign memfont[5944] = 1'd0;
    assign memfont[5945] = 1'd1;
    assign memfont[5946] = 1'd1;
    assign memfont[5947] = 1'd1;
    assign memfont[5948] = 1'd0;
    assign memfont[5949] = 1'd0;
    assign memfont[5950] = 1'd0;
    assign memfont[5951] = 1'd0;
    assign memfont[5952] = 1'd0;
    assign memfont[5953] = 1'd1;
    assign memfont[5954] = 1'd1;
    assign memfont[5955] = 1'd1;
    assign memfont[5956] = 1'd1;
    assign memfont[5957] = 1'd0;
    assign memfont[5958] = 1'd0;
    assign memfont[5959] = 1'd0;
    assign memfont[5960] = 1'd0;
    assign memfont[5961] = 1'd0;
    assign memfont[5962] = 1'd0;
    assign memfont[5963] = 1'd0;
    assign memfont[5964] = 1'd0;
    assign memfont[5965] = 1'd1;
    assign memfont[5966] = 1'd1;
    assign memfont[5967] = 1'd1;
    assign memfont[5968] = 1'd1;
    assign memfont[5969] = 1'd1;
    assign memfont[5970] = 1'd1;
    assign memfont[5971] = 1'd1;
    assign memfont[5972] = 1'd1;
    assign memfont[5973] = 1'd1;
    assign memfont[5974] = 1'd1;
    assign memfont[5975] = 1'd0;
    assign memfont[5976] = 1'd0;
    assign memfont[5977] = 1'd1;
    assign memfont[5978] = 1'd1;
    assign memfont[5979] = 1'd0;
    assign memfont[5980] = 1'd0;
    assign memfont[5981] = 1'd0;
    assign memfont[5982] = 1'd0;
    assign memfont[5983] = 1'd0;
    assign memfont[5984] = 1'd0;
    assign memfont[5985] = 1'd0;
    assign memfont[5986] = 1'd0;
    assign memfont[5987] = 1'd0;
    assign memfont[5988] = 1'd0;
    assign memfont[5989] = 1'd0;
    assign memfont[5990] = 1'd0;
    assign memfont[5991] = 1'd0;
    assign memfont[5992] = 1'd0;
    assign memfont[5993] = 1'd1;
    assign memfont[5994] = 1'd1;
    assign memfont[5995] = 1'd0;
    assign memfont[5996] = 1'd0;
    assign memfont[5997] = 1'd1;
    assign memfont[5998] = 1'd1;
    assign memfont[5999] = 1'd0;
    assign memfont[6000] = 1'd0;
    assign memfont[6001] = 1'd1;
    assign memfont[6002] = 1'd1;
    assign memfont[6003] = 1'd0;
    assign memfont[6004] = 1'd0;
    assign memfont[6005] = 1'd0;
    assign memfont[6006] = 1'd0;
    assign memfont[6007] = 1'd0;
    assign memfont[6008] = 1'd0;
    assign memfont[6009] = 1'd1;
    assign memfont[6010] = 1'd1;
    assign memfont[6011] = 1'd0;
    assign memfont[6012] = 1'd0;
    assign memfont[6013] = 1'd0;
    assign memfont[6014] = 1'd0;
    assign memfont[6015] = 1'd0;
    assign memfont[6016] = 1'd0;
    assign memfont[6017] = 1'd1;
    assign memfont[6018] = 1'd1;
    assign memfont[6019] = 1'd0;
    assign memfont[6020] = 1'd0;
    assign memfont[6021] = 1'd0;
    assign memfont[6022] = 1'd0;
    assign memfont[6023] = 1'd0;
    assign memfont[6024] = 1'd0;
    assign memfont[6025] = 1'd0;
    assign memfont[6026] = 1'd0;
    assign memfont[6027] = 1'd0;
    assign memfont[6028] = 1'd1;
    assign memfont[6029] = 1'd1;
    assign memfont[6030] = 1'd1;
    assign memfont[6031] = 1'd0;
    assign memfont[6032] = 1'd0;
    assign memfont[6033] = 1'd0;
    assign memfont[6034] = 1'd0;
    assign memfont[6035] = 1'd0;
    assign memfont[6036] = 1'd0;
    assign memfont[6037] = 1'd1;
    assign memfont[6038] = 1'd1;
    assign memfont[6039] = 1'd0;
    assign memfont[6040] = 1'd0;
    assign memfont[6041] = 1'd0;
    assign memfont[6042] = 1'd0;
    assign memfont[6043] = 1'd0;
    assign memfont[6044] = 1'd0;
    assign memfont[6045] = 1'd1;
    assign memfont[6046] = 1'd1;
    assign memfont[6047] = 1'd0;
    assign memfont[6048] = 1'd0;
    assign memfont[6049] = 1'd1;
    assign memfont[6050] = 1'd1;
    assign memfont[6051] = 1'd1;
    assign memfont[6052] = 1'd1;
    assign memfont[6053] = 1'd1;
    assign memfont[6054] = 1'd1;
    assign memfont[6055] = 1'd1;
    assign memfont[6056] = 1'd1;
    assign memfont[6057] = 1'd1;
    assign memfont[6058] = 1'd1;
    assign memfont[6059] = 1'd0;
    assign memfont[6060] = 1'd0;
    assign memfont[6061] = 1'd1;
    assign memfont[6062] = 1'd1;
    assign memfont[6063] = 1'd0;
    assign memfont[6064] = 1'd0;
    assign memfont[6065] = 1'd1;
    assign memfont[6066] = 1'd1;
    assign memfont[6067] = 1'd0;
    assign memfont[6068] = 1'd0;
    assign memfont[6069] = 1'd1;
    assign memfont[6070] = 1'd1;
    assign memfont[6071] = 1'd0;
    assign memfont[6072] = 1'd0;
    assign memfont[6073] = 1'd1;
    assign memfont[6074] = 1'd1;
    assign memfont[6075] = 1'd0;
    assign memfont[6076] = 1'd0;
    assign memfont[6077] = 1'd0;
    assign memfont[6078] = 1'd0;
    assign memfont[6079] = 1'd0;
    assign memfont[6080] = 1'd1;
    assign memfont[6081] = 1'd1;
    assign memfont[6082] = 1'd1;
    assign memfont[6083] = 1'd0;
    assign memfont[6084] = 1'd0;
    assign memfont[6085] = 1'd0;
    assign memfont[6086] = 1'd0;
    assign memfont[6087] = 1'd0;
    assign memfont[6088] = 1'd1;
    assign memfont[6089] = 1'd1;
    assign memfont[6090] = 1'd1;
    assign memfont[6091] = 1'd0;
    assign memfont[6092] = 1'd0;
    assign memfont[6093] = 1'd0;
    assign memfont[6094] = 1'd0;
    assign memfont[6095] = 1'd0;
    assign memfont[6096] = 1'd0;
    assign memfont[6097] = 1'd1;
    assign memfont[6098] = 1'd1;
    assign memfont[6099] = 1'd0;
    assign memfont[6100] = 1'd0;
    assign memfont[6101] = 1'd0;
    assign memfont[6102] = 1'd0;
    assign memfont[6103] = 1'd0;
    assign memfont[6104] = 1'd0;
    assign memfont[6105] = 1'd0;
    assign memfont[6106] = 1'd0;
    assign memfont[6107] = 1'd0;
    assign memfont[6108] = 1'd0;
    assign memfont[6109] = 1'd0;
    assign memfont[6110] = 1'd0;
    assign memfont[6111] = 1'd0;
    assign memfont[6112] = 1'd1;
    assign memfont[6113] = 1'd1;
    assign memfont[6114] = 1'd1;
    assign memfont[6115] = 1'd0;
    assign memfont[6116] = 1'd1;
    assign memfont[6117] = 1'd1;
    assign memfont[6118] = 1'd0;
    assign memfont[6119] = 1'd0;
    assign memfont[6120] = 1'd0;
    assign memfont[6121] = 1'd1;
    assign memfont[6122] = 1'd1;
    assign memfont[6123] = 1'd0;
    assign memfont[6124] = 1'd0;
    assign memfont[6125] = 1'd0;
    assign memfont[6126] = 1'd0;
    assign memfont[6127] = 1'd0;
    assign memfont[6128] = 1'd0;
    assign memfont[6129] = 1'd1;
    assign memfont[6130] = 1'd1;
    assign memfont[6131] = 1'd0;
    assign memfont[6132] = 1'd0;
    assign memfont[6133] = 1'd0;
    assign memfont[6134] = 1'd0;
    assign memfont[6135] = 1'd0;
    assign memfont[6136] = 1'd1;
    assign memfont[6137] = 1'd1;
    assign memfont[6138] = 1'd1;
    assign memfont[6139] = 1'd1;
    assign memfont[6140] = 1'd0;
    assign memfont[6141] = 1'd0;
    assign memfont[6142] = 1'd0;
    assign memfont[6143] = 1'd0;
    assign memfont[6144] = 1'd0;
    assign memfont[6145] = 1'd0;
    assign memfont[6146] = 1'd0;
    assign memfont[6147] = 1'd0;
    assign memfont[6148] = 1'd0;
    assign memfont[6149] = 1'd1;
    assign memfont[6150] = 1'd1;
    assign memfont[6151] = 1'd0;
    assign memfont[6152] = 1'd0;
    assign memfont[6153] = 1'd0;
    assign memfont[6154] = 1'd0;
    assign memfont[6155] = 1'd0;
    assign memfont[6156] = 1'd0;
    assign memfont[6157] = 1'd0;
    assign memfont[6158] = 1'd0;
    assign memfont[6159] = 1'd0;
    assign memfont[6160] = 1'd1;
    assign memfont[6161] = 1'd1;
    assign memfont[6162] = 1'd1;
    assign memfont[6163] = 1'd1;
    assign memfont[6164] = 1'd0;
    assign memfont[6165] = 1'd0;
    assign memfont[6166] = 1'd0;
    assign memfont[6167] = 1'd0;
    assign memfont[6168] = 1'd0;
    assign memfont[6169] = 1'd0;
    assign memfont[6170] = 1'd0;
    assign memfont[6171] = 1'd0;
    assign memfont[6172] = 1'd0;
    assign memfont[6173] = 1'd1;
    assign memfont[6174] = 1'd1;
    assign memfont[6175] = 1'd0;
    assign memfont[6176] = 1'd0;
    assign memfont[6177] = 1'd0;
    assign memfont[6178] = 1'd0;
    assign memfont[6179] = 1'd0;
    assign memfont[6180] = 1'd0;
    assign memfont[6181] = 1'd0;
    assign memfont[6182] = 1'd1;
    assign memfont[6183] = 1'd1;
    assign memfont[6184] = 1'd0;
    assign memfont[6185] = 1'd0;
    assign memfont[6186] = 1'd0;
    assign memfont[6187] = 1'd0;
    assign memfont[6188] = 1'd1;
    assign memfont[6189] = 1'd0;
    assign memfont[6190] = 1'd0;
    assign memfont[6191] = 1'd0;
    assign memfont[6192] = 1'd1;
    assign memfont[6193] = 1'd1;
    assign memfont[6194] = 1'd1;
    assign memfont[6195] = 1'd0;
    assign memfont[6196] = 1'd0;
    assign memfont[6197] = 1'd0;
    assign memfont[6198] = 1'd0;
    assign memfont[6199] = 1'd0;
    assign memfont[6200] = 1'd0;
    assign memfont[6201] = 1'd1;
    assign memfont[6202] = 1'd1;
    assign memfont[6203] = 1'd0;
    assign memfont[6204] = 1'd0;
    assign memfont[6205] = 1'd0;
    assign memfont[6206] = 1'd0;
    assign memfont[6207] = 1'd0;
    assign memfont[6208] = 1'd0;
    assign memfont[6209] = 1'd1;
    assign memfont[6210] = 1'd1;
    assign memfont[6211] = 1'd0;
    assign memfont[6212] = 1'd0;
    assign memfont[6213] = 1'd0;
    assign memfont[6214] = 1'd0;
    assign memfont[6215] = 1'd0;
    assign memfont[6216] = 1'd0;
    assign memfont[6217] = 1'd1;
    assign memfont[6218] = 1'd1;
    assign memfont[6219] = 1'd1;
    assign memfont[6220] = 1'd1;
    assign memfont[6221] = 1'd1;
    assign memfont[6222] = 1'd1;
    assign memfont[6223] = 1'd1;
    assign memfont[6224] = 1'd1;
    assign memfont[6225] = 1'd1;
    assign memfont[6226] = 1'd1;
    assign memfont[6227] = 1'd0;
    assign memfont[6228] = 1'd0;
    assign memfont[6229] = 1'd0;
    assign memfont[6230] = 1'd0;
    assign memfont[6231] = 1'd0;
    assign memfont[6232] = 1'd1;
    assign memfont[6233] = 1'd1;
    assign memfont[6234] = 1'd1;
    assign memfont[6235] = 1'd0;
    assign memfont[6236] = 1'd0;
    assign memfont[6237] = 1'd0;
    assign memfont[6238] = 1'd0;
    assign memfont[6239] = 1'd0;
    assign memfont[6240] = 1'd0;
    assign memfont[6241] = 1'd0;
    assign memfont[6242] = 1'd0;
    assign memfont[6243] = 1'd0;
    assign memfont[6244] = 1'd0;
    assign memfont[6245] = 1'd0;
    assign memfont[6246] = 1'd0;
    assign memfont[6247] = 1'd0;
    assign memfont[6248] = 1'd0;
    assign memfont[6249] = 1'd0;
    assign memfont[6250] = 1'd0;
    assign memfont[6251] = 1'd0;
    assign memfont[6252] = 1'd0;
    assign memfont[6253] = 1'd0;
    assign memfont[6254] = 1'd0;
    assign memfont[6255] = 1'd0;
    assign memfont[6256] = 1'd0;
    assign memfont[6257] = 1'd0;
    assign memfont[6258] = 1'd0;
    assign memfont[6259] = 1'd0;
    assign memfont[6260] = 1'd0;
    assign memfont[6261] = 1'd0;
    assign memfont[6262] = 1'd0;
    assign memfont[6263] = 1'd0;


endmodule
