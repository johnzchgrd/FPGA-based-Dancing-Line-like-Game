module hat_rom (
    input clk,
	output reg [5:0] dout,
	input [11:0] addr
    );
	
	wire [5:0] memory [4095:0];

	always @(posedge clk) begin
        dout = memory[addr[11:0]];
    end
    
    assign memory[0   ] = 6'd32;
    assign memory[1   ] = 6'd31;
    assign memory[2   ] = 6'd32;
    assign memory[3   ] = 6'd32;
    assign memory[4   ] = 6'd32;
    assign memory[5   ] = 6'd30;
    assign memory[6   ] = 6'd25;
    assign memory[7   ] = 6'd22;
    assign memory[8   ] = 6'd25;
    assign memory[9   ] = 6'd29;
    assign memory[10  ] = 6'd30;
    assign memory[11  ] = 6'd30;
    assign memory[12  ] = 6'd30;
    assign memory[13  ] = 6'd30;
    assign memory[14  ] = 6'd30;
    assign memory[15  ] = 6'd30;
    assign memory[16  ] = 6'd30;
    assign memory[17  ] = 6'd31;
    assign memory[18  ] = 6'd36;
    assign memory[19  ] = 6'd37;
    assign memory[20  ] = 6'd37;
    assign memory[21  ] = 6'd40;
    assign memory[22  ] = 6'd41;
    assign memory[23  ] = 6'd39;
    assign memory[24  ] = 6'd37;
    assign memory[25  ] = 6'd37;
    assign memory[26  ] = 6'd35;
    assign memory[27  ] = 6'd30;
    assign memory[28  ] = 6'd32;
    assign memory[29  ] = 6'd23;
    assign memory[30  ] = 6'd8 ;
    assign memory[31  ] = 6'd3 ;
    assign memory[32  ] = 6'd12;
    assign memory[33  ] = 6'd28;
    assign memory[34  ] = 6'd31;
    assign memory[35  ] = 6'd29;
    assign memory[36  ] = 6'd30;
    assign memory[37  ] = 6'd30;
    assign memory[38  ] = 6'd30;
    assign memory[39  ] = 6'd30;
    assign memory[40  ] = 6'd30;
    assign memory[41  ] = 6'd30;
    assign memory[42  ] = 6'd30;
    assign memory[43  ] = 6'd30;
    assign memory[44  ] = 6'd30;
    assign memory[45  ] = 6'd30;
    assign memory[46  ] = 6'd30;
    assign memory[47  ] = 6'd30;
    assign memory[48  ] = 6'd31;
    assign memory[49  ] = 6'd29;
    assign memory[50  ] = 6'd30;
    assign memory[51  ] = 6'd30;
    assign memory[52  ] = 6'd30;
    assign memory[53  ] = 6'd30;
    assign memory[54  ] = 6'd30;
    assign memory[55  ] = 6'd30;
    assign memory[56  ] = 6'd30;
    assign memory[57  ] = 6'd30;
    assign memory[58  ] = 6'd30;
    assign memory[59  ] = 6'd30;
    assign memory[60  ] = 6'd30;
    assign memory[61  ] = 6'd30;
    assign memory[62  ] = 6'd30;
    assign memory[63  ] = 6'd30;
    assign memory[64  ] = 6'd30;
    assign memory[65  ] = 6'd30;
    assign memory[66  ] = 6'd30;
    assign memory[67  ] = 6'd30;
    assign memory[68  ] = 6'd30;
    assign memory[69  ] = 6'd29;
    assign memory[70  ] = 6'd30;
    assign memory[71  ] = 6'd30;
    assign memory[72  ] = 6'd30;
    assign memory[73  ] = 6'd30;
    assign memory[74  ] = 6'd30;
    assign memory[75  ] = 6'd30;
    assign memory[76  ] = 6'd30;
    assign memory[77  ] = 6'd30;
    assign memory[78  ] = 6'd30;
    assign memory[79  ] = 6'd30;
    assign memory[80  ] = 6'd30;
    assign memory[81  ] = 6'd30;
    assign memory[82  ] = 6'd31;
    assign memory[83  ] = 6'd27;
    assign memory[84  ] = 6'd14;
    assign memory[85  ] = 6'd12;
    assign memory[86  ] = 6'd12;
    assign memory[87  ] = 6'd7 ;
    assign memory[88  ] = 6'd4 ;
    assign memory[89  ] = 6'd13;
    assign memory[90  ] = 6'd33;
    assign memory[91  ] = 6'd40;
    assign memory[92  ] = 6'd33;
    assign memory[93  ] = 6'd22;
    assign memory[94  ] = 6'd18;
    assign memory[95  ] = 6'd24;
    assign memory[96  ] = 6'd38;
    assign memory[97  ] = 6'd41;
    assign memory[98  ] = 6'd41;
    assign memory[99  ] = 6'd43;
    assign memory[100 ] = 6'd45;
    assign memory[101 ] = 6'd42;
    assign memory[102 ] = 6'd34;
    assign memory[103 ] = 6'd32;
    assign memory[104 ] = 6'd36;
    assign memory[105 ] = 6'd46;
    assign memory[106 ] = 6'd47;
    assign memory[107 ] = 6'd49;
    assign memory[108 ] = 6'd56;
    assign memory[109 ] = 6'd58;
    assign memory[110 ] = 6'd57;
    assign memory[111 ] = 6'd57;
    assign memory[112 ] = 6'd60;
    assign memory[113 ] = 6'd49;
    assign memory[114 ] = 6'd20;
    assign memory[115 ] = 6'd8 ;
    assign memory[116 ] = 6'd20;
    assign memory[117 ] = 6'd38;
    assign memory[118 ] = 6'd47;
    assign memory[119 ] = 6'd40;
    assign memory[120 ] = 6'd33;
    assign memory[121 ] = 6'd27;
    assign memory[122 ] = 6'd35;
    assign memory[123 ] = 6'd50;
    assign memory[124 ] = 6'd58;
    assign memory[125 ] = 6'd45;
    assign memory[126 ] = 6'd13;
    assign memory[127 ] = 6'd0 ;
    assign memory[128 ] = 6'd17;
    assign memory[129 ] = 6'd50;
    assign memory[130 ] = 6'd62;
    assign memory[131 ] = 6'd52;
    assign memory[132 ] = 6'd36;
    assign memory[133 ] = 6'd34;
    assign memory[134 ] = 6'd29;
    assign memory[135 ] = 6'd10;
    assign memory[136 ] = 6'd3 ;
    assign memory[137 ] = 6'd13;
    assign memory[138 ] = 6'd36;
    assign memory[139 ] = 6'd42;
    assign memory[140 ] = 6'd40;
    assign memory[141 ] = 6'd40;
    assign memory[142 ] = 6'd42;
    assign memory[143 ] = 6'd35;
    assign memory[144 ] = 6'd15;
    assign memory[145 ] = 6'd6 ;
    assign memory[146 ] = 6'd15;
    assign memory[147 ] = 6'd35;
    assign memory[148 ] = 6'd42;
    assign memory[149 ] = 6'd38;
    assign memory[150 ] = 6'd31;
    assign memory[151 ] = 6'd29;
    assign memory[152 ] = 6'd30;
    assign memory[153 ] = 6'd30;
    assign memory[154 ] = 6'd31;
    assign memory[155 ] = 6'd27;
    assign memory[156 ] = 6'd16;
    assign memory[157 ] = 6'd11;
    assign memory[158 ] = 6'd14;
    assign memory[159 ] = 6'd19;
    assign memory[160 ] = 6'd20;
    assign memory[161 ] = 6'd20;
    assign memory[162 ] = 6'd23;
    assign memory[163 ] = 6'd22;
    assign memory[164 ] = 6'd26;
    assign memory[165 ] = 6'd37;
    assign memory[166 ] = 6'd44;
    assign memory[167 ] = 6'd34;
    assign memory[168 ] = 6'd12;
    assign memory[169 ] = 6'd3 ;
    assign memory[170 ] = 6'd9 ;
    assign memory[171 ] = 6'd15;
    assign memory[172 ] = 6'd18;
    assign memory[173 ] = 6'd15;
    assign memory[174 ] = 6'd11;
    assign memory[175 ] = 6'd10;
    assign memory[176 ] = 6'd9 ;
    assign memory[177 ] = 6'd11;
    assign memory[178 ] = 6'd6 ;
    assign memory[179 ] = 6'd18;
    assign memory[180 ] = 6'd48;
    assign memory[181 ] = 6'd63;
    assign memory[182 ] = 6'd51;
    assign memory[183 ] = 6'd27;
    assign memory[184 ] = 6'd17;
    assign memory[185 ] = 6'd22;
    assign memory[186 ] = 6'd29;
    assign memory[187 ] = 6'd31;
    assign memory[188 ] = 6'd30;
    assign memory[189 ] = 6'd30;
    assign memory[190 ] = 6'd31;
    assign memory[191 ] = 6'd29;
    assign memory[192 ] = 6'd28;
    assign memory[193 ] = 6'd24;
    assign memory[194 ] = 6'd31;
    assign memory[195 ] = 6'd51;
    assign memory[196 ] = 6'd61;
    assign memory[197 ] = 6'd54;
    assign memory[198 ] = 6'd39;
    assign memory[199 ] = 6'd31;
    assign memory[200 ] = 6'd37;
    assign memory[201 ] = 6'd52;
    assign memory[202 ] = 6'd62;
    assign memory[203 ] = 6'd52;
    assign memory[204 ] = 6'd31;
    assign memory[205 ] = 6'd20;
    assign memory[206 ] = 6'd26;
    assign memory[207 ] = 6'd37;
    assign memory[208 ] = 6'd41;
    assign memory[209 ] = 6'd41;
    assign memory[210 ] = 6'd46;
    assign memory[211 ] = 6'd48;
    assign memory[212 ] = 6'd47;
    assign memory[213 ] = 6'd49;
    assign memory[214 ] = 6'd52;
    assign memory[215 ] = 6'd48;
    assign memory[216 ] = 6'd32;
    assign memory[217 ] = 6'd24;
    assign memory[218 ] = 6'd29;
    assign memory[219 ] = 6'd32;
    assign memory[220 ] = 6'd34;
    assign memory[221 ] = 6'd32;
    assign memory[222 ] = 6'd23;
    assign memory[223 ] = 6'd18;
    assign memory[224 ] = 6'd24;
    assign memory[225 ] = 6'd46;
    assign memory[226 ] = 6'd59;
    assign memory[227 ] = 6'd47;
    assign memory[228 ] = 6'd17;
    assign memory[229 ] = 6'd1 ;
    assign memory[230 ] = 6'd10;
    assign memory[231 ] = 6'd25;
    assign memory[232 ] = 6'd32;
    assign memory[233 ] = 6'd30;
    assign memory[234 ] = 6'd30;
    assign memory[235 ] = 6'd30;
    assign memory[236 ] = 6'd30;
    assign memory[237 ] = 6'd24;
    assign memory[238 ] = 6'd23;
    assign memory[239 ] = 6'd23;
    assign memory[240 ] = 6'd27;
    assign memory[241 ] = 6'd25;
    assign memory[242 ] = 6'd28;
    assign memory[243 ] = 6'd41;
    assign memory[244 ] = 6'd46;
    assign memory[245 ] = 6'd42;
    assign memory[246 ] = 6'd33;
    assign memory[247 ] = 6'd30;
    assign memory[248 ] = 6'd29;
    assign memory[249 ] = 6'd23;
    assign memory[250 ] = 6'd18;
    assign memory[251 ] = 6'd23;
    assign memory[252 ] = 6'd38;
    assign memory[253 ] = 6'd47;
    assign memory[254 ] = 6'd41;
    assign memory[255 ] = 6'd26;
    assign memory[256 ] = 6'd17;
    assign memory[257 ] = 6'd22;
    assign memory[258 ] = 6'd35;
    assign memory[259 ] = 6'd42;
    assign memory[260 ] = 6'd39;
    assign memory[261 ] = 6'd35;
    assign memory[262 ] = 6'd32;
    assign memory[263 ] = 6'd36;
    assign memory[264 ] = 6'd50;
    assign memory[265 ] = 6'd62;
    assign memory[266 ] = 6'd53;
    assign memory[267 ] = 6'd24;
    assign memory[268 ] = 6'd9 ;
    assign memory[269 ] = 6'd15;
    assign memory[270 ] = 6'd26;
    assign memory[271 ] = 6'd30;
    assign memory[272 ] = 6'd32;
    assign memory[273 ] = 6'd50;
    assign memory[274 ] = 6'd59;
    assign memory[275 ] = 6'd57;
    assign memory[276 ] = 6'd51;
    assign memory[277 ] = 6'd52;
    assign memory[278 ] = 6'd47;
    assign memory[279 ] = 6'd28;
    assign memory[280 ] = 6'd16;
    assign memory[281 ] = 6'd23;
    assign memory[282 ] = 6'd48;
    assign memory[283 ] = 6'd62;
    assign memory[284 ] = 6'd54;
    assign memory[285 ] = 6'd27;
    assign memory[286 ] = 6'd12;
    assign memory[287 ] = 6'd20;
    assign memory[288 ] = 6'd44;
    assign memory[289 ] = 6'd58;
    assign memory[290 ] = 6'd51;
    assign memory[291 ] = 6'd39;
    assign memory[292 ] = 6'd32;
    assign memory[293 ] = 6'd34;
    assign memory[294 ] = 6'd31;
    assign memory[295 ] = 6'd30;
    assign memory[296 ] = 6'd31;
    assign memory[297 ] = 6'd35;
    assign memory[298 ] = 6'd37;
    assign memory[299 ] = 6'd37;
    assign memory[300 ] = 6'd41;
    assign memory[301 ] = 6'd46;
    assign memory[302 ] = 6'd40;
    assign memory[303 ] = 6'd22;
    assign memory[304 ] = 6'd9 ;
    assign memory[305 ] = 6'd16;
    assign memory[306 ] = 6'd40;
    assign memory[307 ] = 6'd54;
    assign memory[308 ] = 6'd48;
    assign memory[309 ] = 6'd23;
    assign memory[310 ] = 6'd11;
    assign memory[311 ] = 6'd14;
    assign memory[312 ] = 6'd23;
    assign memory[313 ] = 6'd26;
    assign memory[314 ] = 6'd28;
    assign memory[315 ] = 6'd45;
    assign memory[316 ] = 6'd58;
    assign memory[317 ] = 6'd50;
    assign memory[318 ] = 6'd20;
    assign memory[319 ] = 6'd1 ;
    assign memory[320 ] = 6'd8 ;
    assign memory[321 ] = 6'd29;
    assign memory[322 ] = 6'd39;
    assign memory[323 ] = 6'd36;
    assign memory[324 ] = 6'd32;
    assign memory[325 ] = 6'd30;
    assign memory[326 ] = 6'd30;
    assign memory[327 ] = 6'd18;
    assign memory[328 ] = 6'd11;
    assign memory[329 ] = 6'd14;
    assign memory[330 ] = 6'd20;
    assign memory[331 ] = 6'd24;
    assign memory[332 ] = 6'd23;
    assign memory[333 ] = 6'd21;
    assign memory[334 ] = 6'd20;
    assign memory[335 ] = 6'd20;
    assign memory[336 ] = 6'd13;
    assign memory[337 ] = 6'd7 ;
    assign memory[338 ] = 6'd11;
    assign memory[339 ] = 6'd35;
    assign memory[340 ] = 6'd52;
    assign memory[341 ] = 6'd45;
    assign memory[342 ] = 6'd20;
    assign memory[343 ] = 6'd3 ;
    assign memory[344 ] = 6'd8 ;
    assign memory[345 ] = 6'd25;
    assign memory[346 ] = 6'd35;
    assign memory[347 ] = 6'd34;
    assign memory[348 ] = 6'd31;
    assign memory[349 ] = 6'd29;
    assign memory[350 ] = 6'd31;
    assign memory[351 ] = 6'd34;
    assign memory[352 ] = 6'd38;
    assign memory[353 ] = 6'd36;
    assign memory[354 ] = 6'd29;
    assign memory[355 ] = 6'd22;
    assign memory[356 ] = 6'd24;
    assign memory[357 ] = 6'd33;
    assign memory[358 ] = 6'd38;
    assign memory[359 ] = 6'd37;
    assign memory[360 ] = 6'd32;
    assign memory[361 ] = 6'd30;
    assign memory[362 ] = 6'd30;
    assign memory[363 ] = 6'd38;
    assign memory[364 ] = 6'd40;
    assign memory[365 ] = 6'd41;
    assign memory[366 ] = 6'd42;
    assign memory[367 ] = 6'd46;
    assign memory[368 ] = 6'd43;
    assign memory[369 ] = 6'd19;
    assign memory[370 ] = 6'd3 ;
    assign memory[371 ] = 6'd8 ;
    assign memory[372 ] = 6'd39;
    assign memory[373 ] = 6'd57;
    assign memory[374 ] = 6'd53;
    assign memory[375 ] = 6'd43;
    assign memory[376 ] = 6'd35;
    assign memory[377 ] = 6'd38;
    assign memory[378 ] = 6'd41;
    assign memory[379 ] = 6'd46;
    assign memory[380 ] = 6'd43;
    assign memory[381 ] = 6'd26;
    assign memory[382 ] = 6'd14;
    assign memory[383 ] = 6'd17;
    assign memory[384 ] = 6'd29;
    assign memory[385 ] = 6'd34;
    assign memory[386 ] = 6'd34;
    assign memory[387 ] = 6'd35;
    assign memory[388 ] = 6'd38;
    assign memory[389 ] = 6'd36;
    assign memory[390 ] = 6'd29;
    assign memory[391 ] = 6'd22;
    assign memory[392 ] = 6'd24;
    assign memory[393 ] = 6'd36;
    assign memory[394 ] = 6'd45;
    assign memory[395 ] = 6'd43;
    assign memory[396 ] = 6'd43;
    assign memory[397 ] = 6'd45;
    assign memory[398 ] = 6'd43;
    assign memory[399 ] = 6'd29;
    assign memory[400 ] = 6'd17;
    assign memory[401 ] = 6'd21;
    assign memory[402 ] = 6'd29;
    assign memory[403 ] = 6'd35;
    assign memory[404 ] = 6'd33;
    assign memory[405 ] = 6'd27;
    assign memory[406 ] = 6'd22;
    assign memory[407 ] = 6'd23;
    assign memory[408 ] = 6'd33;
    assign memory[409 ] = 6'd38;
    assign memory[410 ] = 6'd37;
    assign memory[411 ] = 6'd34;
    assign memory[412 ] = 6'd33;
    assign memory[413 ] = 6'd33;
    assign memory[414 ] = 6'd38;
    assign memory[415 ] = 6'd41;
    assign memory[416 ] = 6'd40;
    assign memory[417 ] = 6'd37;
    assign memory[418 ] = 6'd37;
    assign memory[419 ] = 6'd37;
    assign memory[420 ] = 6'd25;
    assign memory[421 ] = 6'd15;
    assign memory[422 ] = 6'd17;
    assign memory[423 ] = 6'd38;
    assign memory[424 ] = 6'd53;
    assign memory[425 ] = 6'd49;
    assign memory[426 ] = 6'd40;
    assign memory[427 ] = 6'd32;
    assign memory[428 ] = 6'd34;
    assign memory[429 ] = 6'd42;
    assign memory[430 ] = 6'd49;
    assign memory[431 ] = 6'd47;
    assign memory[432 ] = 6'd36;
    assign memory[433 ] = 6'd30;
    assign memory[434 ] = 6'd29;
    assign memory[435 ] = 6'd31;
    assign memory[436 ] = 6'd29;
    assign memory[437 ] = 6'd31;
    assign memory[438 ] = 6'd38;
    assign memory[439 ] = 6'd45;
    assign memory[440 ] = 6'd44;
    assign memory[441 ] = 6'd38;
    assign memory[442 ] = 6'd32;
    assign memory[443 ] = 6'd33;
    assign memory[444 ] = 6'd41;
    assign memory[445 ] = 6'd48;
    assign memory[446 ] = 6'd47;
    assign memory[447 ] = 6'd32;
    assign memory[448 ] = 6'd22;
    assign memory[449 ] = 6'd23;
    assign memory[450 ] = 6'd29;
    assign memory[451 ] = 6'd35;
    assign memory[452 ] = 6'd33;
    assign memory[453 ] = 6'd29;
    assign memory[454 ] = 6'd25;
    assign memory[455 ] = 6'd27;
    assign memory[456 ] = 6'd38;
    assign memory[457 ] = 6'd49;
    assign memory[458 ] = 6'd47;
    assign memory[459 ] = 6'd36;
    assign memory[460 ] = 6'd30;
    assign memory[461 ] = 6'd30;
    assign memory[462 ] = 6'd26;
    assign memory[463 ] = 6'd22;
    assign memory[464 ] = 6'd24;
    assign memory[465 ] = 6'd26;
    assign memory[466 ] = 6'd31;
    assign memory[467 ] = 6'd30;
    assign memory[468 ] = 6'd17;
    assign memory[469 ] = 6'd4 ;
    assign memory[470 ] = 6'd5 ;
    assign memory[471 ] = 6'd24;
    assign memory[472 ] = 6'd38;
    assign memory[473 ] = 6'd37;
    assign memory[474 ] = 6'd31;
    assign memory[475 ] = 6'd26;
    assign memory[476 ] = 6'd27;
    assign memory[477 ] = 6'd23;
    assign memory[478 ] = 6'd19;
    assign memory[479 ] = 6'd20;
    assign memory[480 ] = 6'd27;
    assign memory[481 ] = 6'd34;
    assign memory[482 ] = 6'd34;
    assign memory[483 ] = 6'd27;
    assign memory[484 ] = 6'd23;
    assign memory[485 ] = 6'd23;
    assign memory[486 ] = 6'd35;
    assign memory[487 ] = 6'd45;
    assign memory[488 ] = 6'd44;
    assign memory[489 ] = 6'd38;
    assign memory[490 ] = 6'd33;
    assign memory[491 ] = 6'd34;
    assign memory[492 ] = 6'd29;
    assign memory[493 ] = 6'd23;
    assign memory[494 ] = 6'd23;
    assign memory[495 ] = 6'd31;
    assign memory[496 ] = 6'd38;
    assign memory[497 ] = 6'd37;
    assign memory[498 ] = 6'd39;
    assign memory[499 ] = 6'd40;
    assign memory[500 ] = 6'd41;
    assign memory[501 ] = 6'd36;
    assign memory[502 ] = 6'd34;
    assign memory[503 ] = 6'd33;
    assign memory[504 ] = 6'd29;
    assign memory[505 ] = 6'd22;
    assign memory[506 ] = 6'd23;
    assign memory[507 ] = 6'd33;
    assign memory[508 ] = 6'd41;
    assign memory[509 ] = 6'd41;
    assign memory[510 ] = 6'd28;
    assign memory[511 ] = 6'd18;
    assign memory[512 ] = 6'd19;
    assign memory[513 ] = 6'd31;
    assign memory[514 ] = 6'd42;
    assign memory[515 ] = 6'd40;
    assign memory[516 ] = 6'd33;
    assign memory[517 ] = 6'd26;
    assign memory[518 ] = 6'd26;
    assign memory[519 ] = 6'd34;
    assign memory[520 ] = 6'd40;
    assign memory[521 ] = 6'd40;
    assign memory[522 ] = 6'd34;
    assign memory[523 ] = 6'd30;
    assign memory[524 ] = 6'd29;
    assign memory[525 ] = 6'd29;
    assign memory[526 ] = 6'd25;
    assign memory[527 ] = 6'd26;
    assign memory[528 ] = 6'd35;
    assign memory[529 ] = 6'd45;
    assign memory[530 ] = 6'd44;
    assign memory[531 ] = 6'd25;
    assign memory[532 ] = 6'd9 ;
    assign memory[533 ] = 6'd8 ;
    assign memory[534 ] = 6'd19;
    assign memory[535 ] = 6'd27;
    assign memory[536 ] = 6'd27;
    assign memory[537 ] = 6'd30;
    assign memory[538 ] = 6'd33;
    assign memory[539 ] = 6'd34;
    assign memory[540 ] = 6'd30;
    assign memory[541 ] = 6'd26;
    assign memory[542 ] = 6'd27;
    assign memory[543 ] = 6'd25;
    assign memory[544 ] = 6'd23;
    assign memory[545 ] = 6'd23;
    assign memory[546 ] = 6'd28;
    assign memory[547 ] = 6'd31;
    assign memory[548 ] = 6'd31;
    assign memory[549 ] = 6'd29;
    assign memory[550 ] = 6'd27;
    assign memory[551 ] = 6'd27;
    assign memory[552 ] = 6'd32;
    assign memory[553 ] = 6'd38;
    assign memory[554 ] = 6'd38;
    assign memory[555 ] = 6'd28;
    assign memory[556 ] = 6'd19;
    assign memory[557 ] = 6'd18;
    assign memory[558 ] = 6'd30;
    assign memory[559 ] = 6'd41;
    assign memory[560 ] = 6'd41;
    assign memory[561 ] = 6'd31;
    assign memory[562 ] = 6'd22;
    assign memory[563 ] = 6'd22;
    assign memory[564 ] = 6'd26;
    assign memory[565 ] = 6'd31;
    assign memory[566 ] = 6'd29;
    assign memory[567 ] = 6'd36;
    assign memory[568 ] = 6'd44;
    assign memory[569 ] = 6'd43;
    assign memory[570 ] = 6'd39;
    assign memory[571 ] = 6'd34;
    assign memory[572 ] = 6'd34;
    assign memory[573 ] = 6'd29;
    assign memory[574 ] = 6'd23;
    assign memory[575 ] = 6'd23;
    assign memory[576 ] = 6'd28;
    assign memory[577 ] = 6'd33;
    assign memory[578 ] = 6'd33;
    assign memory[579 ] = 6'd36;
    assign memory[580 ] = 6'd40;
    assign memory[581 ] = 6'd41;
    assign memory[582 ] = 6'd37;
    assign memory[583 ] = 6'd34;
    assign memory[584 ] = 6'd33;
    assign memory[585 ] = 6'd34;
    assign memory[586 ] = 6'd33;
    assign memory[587 ] = 6'd34;
    assign memory[588 ] = 6'd29;
    assign memory[589 ] = 6'd23;
    assign memory[590 ] = 6'd23;
    assign memory[591 ] = 6'd25;
    assign memory[592 ] = 6'd26;
    assign memory[593 ] = 6'd26;
    assign memory[594 ] = 6'd34;
    assign memory[595 ] = 6'd41;
    assign memory[596 ] = 6'd42;
    assign memory[597 ] = 6'd32;
    assign memory[598 ] = 6'd23;
    assign memory[599 ] = 6'd23;
    assign memory[600 ] = 6'd19;
    assign memory[601 ] = 6'd13;
    assign memory[602 ] = 6'd13;
    assign memory[603 ] = 6'd19;
    assign memory[604 ] = 6'd28;
    assign memory[605 ] = 6'd28;
    assign memory[606 ] = 6'd25;
    assign memory[607 ] = 6'd24;
    assign memory[608 ] = 6'd23;
    assign memory[609 ] = 6'd27;
    assign memory[610 ] = 6'd31;
    assign memory[611 ] = 6'd31;
    assign memory[612 ] = 6'd24;
    assign memory[613 ] = 6'd16;
    assign memory[614 ] = 6'd16;
    assign memory[615 ] = 6'd21;
    assign memory[616 ] = 6'd26;
    assign memory[617 ] = 6'd27;
    assign memory[618 ] = 6'd25;
    assign memory[619 ] = 6'd24;
    assign memory[620 ] = 6'd22;
    assign memory[621 ] = 6'd36;
    assign memory[622 ] = 6'd51;
    assign memory[623 ] = 6'd52;
    assign memory[624 ] = 6'd43;
    assign memory[625 ] = 6'd34;
    assign memory[626 ] = 6'd34;
    assign memory[627 ] = 6'd30;
    assign memory[628 ] = 6'd23;
    assign memory[629 ] = 6'd23;
    assign memory[630 ] = 6'd29;
    assign memory[631 ] = 6'd34;
    assign memory[632 ] = 6'd34;
    assign memory[633 ] = 6'd35;
    assign memory[634 ] = 6'd37;
    assign memory[635 ] = 6'd37;
    assign memory[636 ] = 6'd37;
    assign memory[637 ] = 6'd37;
    assign memory[638 ] = 6'd38;
    assign memory[639 ] = 6'd31;
    assign memory[640 ] = 6'd23;
    assign memory[641 ] = 6'd23;
    assign memory[642 ] = 6'd26;
    assign memory[643 ] = 6'd30;
    assign memory[644 ] = 6'd30;
    assign memory[645 ] = 6'd35;
    assign memory[646 ] = 6'd44;
    assign memory[647 ] = 6'd44;
    assign memory[648 ] = 6'd43;
    assign memory[649 ] = 6'd40;
    assign memory[650 ] = 6'd40;
    assign memory[651 ] = 6'd42;
    assign memory[652 ] = 6'd44;
    assign memory[653 ] = 6'd44;
    assign memory[654 ] = 6'd41;
    assign memory[655 ] = 6'd37;
    assign memory[656 ] = 6'd36;
    assign memory[657 ] = 6'd34;
    assign memory[658 ] = 6'd30;
    assign memory[659 ] = 6'd29;
    assign memory[660 ] = 6'd37;
    assign memory[661 ] = 6'd47;
    assign memory[662 ] = 6'd47;
    assign memory[663 ] = 6'd43;
    assign memory[664 ] = 6'd37;
    assign memory[665 ] = 6'd36;
    assign memory[666 ] = 6'd34;
    assign memory[667 ] = 6'd30;
    assign memory[668 ] = 6'd31;
    assign memory[669 ] = 6'd27;
    assign memory[670 ] = 6'd23;
    assign memory[671 ] = 6'd22;
    assign memory[672 ] = 6'd27;
    assign memory[673 ] = 6'd30;
    assign memory[674 ] = 6'd29;
    assign memory[675 ] = 6'd31;
    assign memory[676 ] = 6'd34;
    assign memory[677 ] = 6'd35;
    assign memory[678 ] = 6'd31;
    assign memory[679 ] = 6'd27;
    assign memory[680 ] = 6'd26;
    assign memory[681 ] = 6'd28;
    assign memory[682 ] = 6'd30;
    assign memory[683 ] = 6'd31;
    assign memory[684 ] = 6'd28;
    assign memory[685 ] = 6'd27;
    assign memory[686 ] = 6'd26;
    assign memory[687 ] = 6'd31;
    assign memory[688 ] = 6'd37;
    assign memory[689 ] = 6'd37;
    assign memory[690 ] = 6'd38;
    assign memory[691 ] = 6'd40;
    assign memory[692 ] = 6'd41;
    assign memory[693 ] = 6'd36;
    assign memory[694 ] = 6'd30;
    assign memory[695 ] = 6'd30;
    assign memory[696 ] = 6'd33;
    assign memory[697 ] = 6'd36;
    assign memory[698 ] = 6'd37;
    assign memory[699 ] = 6'd37;
    assign memory[700 ] = 6'd40;
    assign memory[701 ] = 6'd41;
    assign memory[702 ] = 6'd35;
    assign memory[703 ] = 6'd26;
    assign memory[704 ] = 6'd25;
    assign memory[705 ] = 6'd29;
    assign memory[706 ] = 6'd33;
    assign memory[707 ] = 6'd35;
    assign memory[708 ] = 6'd27;
    assign memory[709 ] = 6'd17;
    assign memory[710 ] = 6'd14;
    assign memory[711 ] = 6'd28;
    assign memory[712 ] = 6'd47;
    assign memory[713 ] = 6'd49;
    assign memory[714 ] = 6'd39;
    assign memory[715 ] = 6'd27;
    assign memory[716 ] = 6'd25;
    assign memory[717 ] = 6'd29;
    assign memory[718 ] = 6'd30;
    assign memory[719 ] = 6'd31;
    assign memory[720 ] = 6'd28;
    assign memory[721 ] = 6'd23;
    assign memory[722 ] = 6'd22;
    assign memory[723 ] = 6'd27;
    assign memory[724 ] = 6'd33;
    assign memory[725 ] = 6'd35;
    assign memory[726 ] = 6'd28;
    assign memory[727 ] = 6'd20;
    assign memory[728 ] = 6'd18;
    assign memory[729 ] = 6'd26;
    assign memory[730 ] = 6'd36;
    assign memory[731 ] = 6'd38;
    assign memory[732 ] = 6'd34;
    assign memory[733 ] = 6'd30;
    assign memory[734 ] = 6'd30;
    assign memory[735 ] = 6'd29;
    assign memory[736 ] = 6'd27;
    assign memory[737 ] = 6'd26;
    assign memory[738 ] = 6'd29;
    assign memory[739 ] = 6'd34;
    assign memory[740 ] = 6'd34;
    assign memory[741 ] = 6'd32;
    assign memory[742 ] = 6'd30;
    assign memory[743 ] = 6'd29;
    assign memory[744 ] = 6'd35;
    assign memory[745 ] = 6'd44;
    assign memory[746 ] = 6'd45;
    assign memory[747 ] = 6'd38;
    assign memory[748 ] = 6'd27;
    assign memory[749 ] = 6'd25;
    assign memory[750 ] = 6'd28;
    assign memory[751 ] = 6'd33;
    assign memory[752 ] = 6'd34;
    assign memory[753 ] = 6'd30;
    assign memory[754 ] = 6'd24;
    assign memory[755 ] = 6'd21;
    assign memory[756 ] = 6'd29;
    assign memory[757 ] = 6'd39;
    assign memory[758 ] = 6'd43;
    assign memory[759 ] = 6'd34;
    assign memory[760 ] = 6'd21;
    assign memory[761 ] = 6'd18;
    assign memory[762 ] = 6'd27;
    assign memory[763 ] = 6'd39;
    assign memory[764 ] = 6'd42;
    assign memory[765 ] = 6'd36;
    assign memory[766 ] = 6'd31;
    assign memory[767 ] = 6'd30;
    assign memory[768 ] = 6'd32;
    assign memory[769 ] = 6'd34;
    assign memory[770 ] = 6'd34;
    assign memory[771 ] = 6'd36;
    assign memory[772 ] = 6'd40;
    assign memory[773 ] = 6'd42;
    assign memory[774 ] = 6'd37;
    assign memory[775 ] = 6'd27;
    assign memory[776 ] = 6'd25;
    assign memory[777 ] = 6'd28;
    assign memory[778 ] = 6'd33;
    assign memory[779 ] = 6'd34;
    assign memory[780 ] = 6'd33;
    assign memory[781 ] = 6'd34;
    assign memory[782 ] = 6'd35;
    assign memory[783 ] = 6'd29;
    assign memory[784 ] = 6'd17;
    assign memory[785 ] = 6'd15;
    assign memory[786 ] = 6'd21;
    assign memory[787 ] = 6'd33;
    assign memory[788 ] = 6'd34;
    assign memory[789 ] = 6'd33;
    assign memory[790 ] = 6'd34;
    assign memory[791 ] = 6'd34;
    assign memory[792 ] = 6'd32;
    assign memory[793 ] = 6'd27;
    assign memory[794 ] = 6'd27;
    assign memory[795 ] = 6'd28;
    assign memory[796 ] = 6'd30;
    assign memory[797 ] = 6'd31;
    assign memory[798 ] = 6'd26;
    assign memory[799 ] = 6'd17;
    assign memory[800 ] = 6'd15;
    assign memory[801 ] = 6'd21;
    assign memory[802 ] = 6'd29;
    assign memory[803 ] = 6'd31;
    assign memory[804 ] = 6'd28;
    assign memory[805 ] = 6'd27;
    assign memory[806 ] = 6'd26;
    assign memory[807 ] = 6'd26;
    assign memory[808 ] = 6'd26;
    assign memory[809 ] = 6'd28;
    assign memory[810 ] = 6'd25;
    assign memory[811 ] = 6'd20;
    assign memory[812 ] = 6'd19;
    assign memory[813 ] = 6'd25;
    assign memory[814 ] = 6'd39;
    assign memory[815 ] = 6'd42;
    assign memory[816 ] = 6'd37;
    assign memory[817 ] = 6'd31;
    assign memory[818 ] = 6'd31;
    assign memory[819 ] = 6'd30;
    assign memory[820 ] = 6'd27;
    assign memory[821 ] = 6'd27;
    assign memory[822 ] = 6'd28;
    assign memory[823 ] = 6'd30;
    assign memory[824 ] = 6'd29;
    assign memory[825 ] = 6'd32;
    assign memory[826 ] = 6'd36;
    assign memory[827 ] = 6'd39;
    assign memory[828 ] = 6'd33;
    assign memory[829 ] = 6'd25;
    assign memory[830 ] = 6'd21;
    assign memory[831 ] = 6'd28;
    assign memory[832 ] = 6'd35;
    assign memory[833 ] = 6'd39;
    assign memory[834 ] = 6'd31;
    assign memory[835 ] = 6'd18;
    assign memory[836 ] = 6'd14;
    assign memory[837 ] = 6'd23;
    assign memory[838 ] = 6'd42;
    assign memory[839 ] = 6'd46;
    assign memory[840 ] = 6'd40;
    assign memory[841 ] = 6'd34;
    assign memory[842 ] = 6'd32;
    assign memory[843 ] = 6'd35;
    assign memory[844 ] = 6'd36;
    assign memory[845 ] = 6'd38;
    assign memory[846 ] = 6'd36;
    assign memory[847 ] = 6'd33;
    assign memory[848 ] = 6'd33;
    assign memory[849 ] = 6'd30;
    assign memory[850 ] = 6'd21;
    assign memory[851 ] = 6'd19;
    assign memory[852 ] = 6'd25;
    assign memory[853 ] = 6'd35;
    assign memory[854 ] = 6'd37;
    assign memory[855 ] = 6'd37;
    assign memory[856 ] = 6'd40;
    assign memory[857 ] = 6'd41;
    assign memory[858 ] = 6'd38;
    assign memory[859 ] = 6'd32;
    assign memory[860 ] = 6'd29;
    assign memory[861 ] = 6'd31;
    assign memory[862 ] = 6'd36;
    assign memory[863 ] = 6'd38;
    assign memory[864 ] = 6'd36;
    assign memory[865 ] = 6'd34;
    assign memory[866 ] = 6'd33;
    assign memory[867 ] = 6'd34;
    assign memory[868 ] = 6'd34;
    assign memory[869 ] = 6'd34;
    assign memory[870 ] = 6'd36;
    assign memory[871 ] = 6'd43;
    assign memory[872 ] = 6'd44;
    assign memory[873 ] = 6'd44;
    assign memory[874 ] = 6'd43;
    assign memory[875 ] = 6'd45;
    assign memory[876 ] = 6'd41;
    assign memory[877 ] = 6'd31;
    assign memory[878 ] = 6'd28;
    assign memory[879 ] = 6'd32;
    assign memory[880 ] = 6'd36;
    assign memory[881 ] = 6'd37;
    assign memory[882 ] = 6'd37;
    assign memory[883 ] = 6'd37;
    assign memory[884 ] = 6'd37;
    assign memory[885 ] = 6'd35;
    assign memory[886 ] = 6'd28;
    assign memory[887 ] = 6'd25;
    assign memory[888 ] = 6'd28;
    assign memory[889 ] = 6'd35;
    assign memory[890 ] = 6'd37;
    assign memory[891 ] = 6'd35;
    assign memory[892 ] = 6'd31;
    assign memory[893 ] = 6'd29;
    assign memory[894 ] = 6'd32;
    assign memory[895 ] = 6'd35;
    assign memory[896 ] = 6'd37;
    assign memory[897 ] = 6'd35;
    assign memory[898 ] = 6'd31;
    assign memory[899 ] = 6'd30;
    assign memory[900 ] = 6'd28;
    assign memory[901 ] = 6'd25;
    assign memory[902 ] = 6'd23;
    assign memory[903 ] = 6'd26;
    assign memory[904 ] = 6'd33;
    assign memory[905 ] = 6'd33;
    assign memory[906 ] = 6'd34;
    assign memory[907 ] = 6'd36;
    assign memory[908 ] = 6'd38;
    assign memory[909 ] = 6'd35;
    assign memory[910 ] = 6'd28;
    assign memory[911 ] = 6'd25;
    assign memory[912 ] = 6'd27;
    assign memory[913 ] = 6'd27;
    assign memory[914 ] = 6'd27;
    assign memory[915 ] = 6'd28;
    assign memory[916 ] = 6'd29;
    assign memory[917 ] = 6'd31;
    assign memory[918 ] = 6'd29;
    assign memory[919 ] = 6'd27;
    assign memory[920 ] = 6'd26;
    assign memory[921 ] = 6'd27;
    assign memory[922 ] = 6'd27;
    assign memory[923 ] = 6'd27;
    assign memory[924 ] = 6'd27;
    assign memory[925 ] = 6'd27;
    assign memory[926 ] = 6'd27;
    assign memory[927 ] = 6'd28;
    assign memory[928 ] = 6'd27;
    assign memory[929 ] = 6'd27;
    assign memory[930 ] = 6'd25;
    assign memory[931 ] = 6'd18;
    assign memory[932 ] = 6'd16;
    assign memory[933 ] = 6'd18;
    assign memory[934 ] = 6'd23;
    assign memory[935 ] = 6'd23;
    assign memory[936 ] = 6'd24;
    assign memory[937 ] = 6'd28;
    assign memory[938 ] = 6'd31;
    assign memory[939 ] = 6'd29;
    assign memory[940 ] = 6'd25;
    assign memory[941 ] = 6'd22;
    assign memory[942 ] = 6'd26;
    assign memory[943 ] = 6'd32;
    assign memory[944 ] = 6'd36;
    assign memory[945 ] = 6'd31;
    assign memory[946 ] = 6'd22;
    assign memory[947 ] = 6'd18;
    assign memory[948 ] = 6'd22;
    assign memory[949 ] = 6'd32;
    assign memory[950 ] = 6'd35;
    assign memory[951 ] = 6'd33;
    assign memory[952 ] = 6'd30;
    assign memory[953 ] = 6'd30;
    assign memory[954 ] = 6'd28;
    assign memory[955 ] = 6'd24;
    assign memory[956 ] = 6'd22;
    assign memory[957 ] = 6'd25;
    assign memory[958 ] = 6'd35;
    assign memory[959 ] = 6'd38;
    assign memory[960 ] = 6'd36;
    assign memory[961 ] = 6'd29;
    assign memory[962 ] = 6'd25;
    assign memory[963 ] = 6'd29;
    assign memory[964 ] = 6'd38;
    assign memory[965 ] = 6'd43;
    assign memory[966 ] = 6'd39;
    assign memory[967 ] = 6'd35;
    assign memory[968 ] = 6'd32;
    assign memory[969 ] = 6'd35;
    assign memory[970 ] = 6'd39;
    assign memory[971 ] = 6'd42;
    assign memory[972 ] = 6'd38;
    assign memory[973 ] = 6'd29;
    assign memory[974 ] = 6'd25;
    assign memory[975 ] = 6'd28;
    assign memory[976 ] = 6'd35;
    assign memory[977 ] = 6'd37;
    assign memory[978 ] = 6'd36;
    assign memory[979 ] = 6'd36;
    assign memory[980 ] = 6'd37;
    assign memory[981 ] = 6'd37;
    assign memory[982 ] = 6'd37;
    assign memory[983 ] = 6'd37;
    assign memory[984 ] = 6'd35;
    assign memory[985 ] = 6'd28;
    assign memory[986 ] = 6'd26;
    assign memory[987 ] = 6'd28;
    assign memory[988 ] = 6'd32;
    assign memory[989 ] = 6'd34;
    assign memory[990 ] = 6'd33;
    assign memory[991 ] = 6'd37;
    assign memory[992 ] = 6'd37;
    assign memory[993 ] = 6'd38;
    assign memory[994 ] = 6'd39;
    assign memory[995 ] = 6'd42;
    assign memory[996 ] = 6'd39;
    assign memory[997 ] = 6'd29;
    assign memory[998 ] = 6'd25;
    assign memory[999 ] = 6'd28;
    assign memory[1000] = 6'd35;
    assign memory[1001] = 6'd38;
    assign memory[1002] = 6'd36;
    assign memory[1003] = 6'd34;
    assign memory[1004] = 6'd34;
    assign memory[1005] = 6'd33;
    assign memory[1006] = 6'd31;
    assign memory[1007] = 6'd29;
    assign memory[1008] = 6'd32;
    assign memory[1009] = 6'd38;
    assign memory[1010] = 6'd42;
    assign memory[1011] = 6'd38;
    assign memory[1012] = 6'd24;
    assign memory[1013] = 6'd18;
    assign memory[1014] = 6'd23;
    assign memory[1015] = 6'd34;
    assign memory[1016] = 6'd38;
    assign memory[1017] = 6'd38;
    assign memory[1018] = 6'd40;
    assign memory[1019] = 6'd42;
    assign memory[1020] = 6'd39;
    assign memory[1021] = 6'd35;
    assign memory[1022] = 6'd34;
    assign memory[1023] = 6'd33;
    assign memory[1024] = 6'd32;
    assign memory[1025] = 6'd29;
    assign memory[1026] = 6'd32;
    assign memory[1027] = 6'd36;
    assign memory[1028] = 6'd38;
    assign memory[1029] = 6'd35;
    assign memory[1030] = 6'd28;
    assign memory[1031] = 6'd25;
    assign memory[1032] = 6'd27;
    assign memory[1033] = 6'd35;
    assign memory[1034] = 6'd39;
    assign memory[1035] = 6'd36;
    assign memory[1036] = 6'd29;
    assign memory[1037] = 6'd26;
    assign memory[1038] = 6'd28;
    assign memory[1039] = 6'd32;
    assign memory[1040] = 6'd34;
    assign memory[1041] = 6'd33;
    assign memory[1042] = 6'd33;
    assign memory[1043] = 6'd33;
    assign memory[1044] = 6'd33;
    assign memory[1045] = 6'd31;
    assign memory[1046] = 6'd30;
    assign memory[1047] = 6'd30;
    assign memory[1048] = 6'd33;
    assign memory[1049] = 6'd34;
    assign memory[1050] = 6'd33;
    assign memory[1051] = 6'd33;
    assign memory[1052] = 6'd33;
    assign memory[1053] = 6'd32;
    assign memory[1054] = 6'd28;
    assign memory[1055] = 6'd26;
    assign memory[1056] = 6'd28;
    assign memory[1057] = 6'd33;
    assign memory[1058] = 6'd34;
    assign memory[1059] = 6'd34;
    assign memory[1060] = 6'd38;
    assign memory[1061] = 6'd41;
    assign memory[1062] = 6'd38;
    assign memory[1063] = 6'd29;
    assign memory[1064] = 6'd26;
    assign memory[1065] = 6'd27;
    assign memory[1066] = 6'd26;
    assign memory[1067] = 6'd27;
    assign memory[1068] = 6'd27;
    assign memory[1069] = 6'd27;
    assign memory[1070] = 6'd26;
    assign memory[1071] = 6'd28;
    assign memory[1072] = 6'd38;
    assign memory[1073] = 6'd45;
    assign memory[1074] = 6'd42;
    assign memory[1075] = 6'd31;
    assign memory[1076] = 6'd26;
    assign memory[1077] = 6'd28;
    assign memory[1078] = 6'd29;
    assign memory[1079] = 6'd31;
    assign memory[1080] = 6'd30;
    assign memory[1081] = 6'd30;
    assign memory[1082] = 6'd31;
    assign memory[1083] = 6'd29;
    assign memory[1084] = 6'd23;
    assign memory[1085] = 6'd18;
    assign memory[1086] = 6'd21;
    assign memory[1087] = 6'd32;
    assign memory[1088] = 6'd38;
    assign memory[1089] = 6'd36;
    assign memory[1090] = 6'd32;
    assign memory[1091] = 6'd29;
    assign memory[1092] = 6'd31;
    assign memory[1093] = 6'd33;
    assign memory[1094] = 6'd35;
    assign memory[1095] = 6'd33;
    assign memory[1096] = 6'd28;
    assign memory[1097] = 6'd26;
    assign memory[1098] = 6'd27;
    assign memory[1099] = 6'd32;
    assign memory[1100] = 6'd34;
    assign memory[1101] = 6'd33;
    assign memory[1102] = 6'd31;
    assign memory[1103] = 6'd29;
    assign memory[1104] = 6'd30;
    assign memory[1105] = 6'd33;
    assign memory[1106] = 6'd35;
    assign memory[1107] = 6'd35;
    assign memory[1108] = 6'd32;
    assign memory[1109] = 6'd30;
    assign memory[1110] = 6'd30;
    assign memory[1111] = 6'd27;
    assign memory[1112] = 6'd26;
    assign memory[1113] = 6'd27;
    assign memory[1114] = 6'd30;
    assign memory[1115] = 6'd31;
    assign memory[1116] = 6'd30;
    assign memory[1117] = 6'd30;
    assign memory[1118] = 6'd31;
    assign memory[1119] = 6'd30;
    assign memory[1120] = 6'd28;
    assign memory[1121] = 6'd26;
    assign memory[1122] = 6'd27;
    assign memory[1123] = 6'd34;
    assign memory[1124] = 6'd38;
    assign memory[1125] = 6'd37;
    assign memory[1126] = 6'd32;
    assign memory[1127] = 6'd29;
    assign memory[1128] = 6'd31;
    assign memory[1129] = 6'd34;
    assign memory[1130] = 6'd38;
    assign memory[1131] = 6'd36;
    assign memory[1132] = 6'd27;
    assign memory[1133] = 6'd22;
    assign memory[1134] = 6'd24;
    assign memory[1135] = 6'd29;
    assign memory[1136] = 6'd31;
    assign memory[1137] = 6'd30;
    assign memory[1138] = 6'd33;
    assign memory[1139] = 6'd34;
    assign memory[1140] = 6'd34;
    assign memory[1141] = 6'd33;
    assign memory[1142] = 6'd33;
    assign memory[1143] = 6'd33;
    assign memory[1144] = 6'd31;
    assign memory[1145] = 6'd30;
    assign memory[1146] = 6'd30;
    assign memory[1147] = 6'd31;
    assign memory[1148] = 6'd30;
    assign memory[1149] = 6'd30;
    assign memory[1150] = 6'd34;
    assign memory[1151] = 6'd38;
    assign memory[1152] = 6'd36;
    assign memory[1153] = 6'd31;
    assign memory[1154] = 6'd26;
    assign memory[1155] = 6'd27;
    assign memory[1156] = 6'd34;
    assign memory[1157] = 6'd38;
    assign memory[1158] = 6'd37;
    assign memory[1159] = 6'd32;
    assign memory[1160] = 6'd29;
    assign memory[1161] = 6'd29;
    assign memory[1162] = 6'd32;
    assign memory[1163] = 6'd34;
    assign memory[1164] = 6'd34;
    assign memory[1165] = 6'd36;
    assign memory[1166] = 6'd37;
    assign memory[1167] = 6'd37;
    assign memory[1168] = 6'd33;
    assign memory[1169] = 6'd30;
    assign memory[1170] = 6'd31;
    assign memory[1171] = 6'd37;
    assign memory[1172] = 6'd41;
    assign memory[1173] = 6'd40;
    assign memory[1174] = 6'd38;
    assign memory[1175] = 6'd37;
    assign memory[1176] = 6'd37;
    assign memory[1177] = 6'd35;
    assign memory[1178] = 6'd34;
    assign memory[1179] = 6'd34;
    assign memory[1180] = 6'd34;
    assign memory[1181] = 6'd33;
    assign memory[1182] = 6'd33;
    assign memory[1183] = 6'd33;
    assign memory[1184] = 6'd33;
    assign memory[1185] = 6'd34;
    assign memory[1186] = 6'd36;
    assign memory[1187] = 6'd37;
    assign memory[1188] = 6'd37;
    assign memory[1189] = 6'd35;
    assign memory[1190] = 6'd33;
    assign memory[1191] = 6'd34;
    assign memory[1192] = 6'd34;
    assign memory[1193] = 6'd34;
    assign memory[1194] = 6'd33;
    assign memory[1195] = 6'd33;
    assign memory[1196] = 6'd33;
    assign memory[1197] = 6'd33;
    assign memory[1198] = 6'd33;
    assign memory[1199] = 6'd33;
    assign memory[1200] = 6'd34;
    assign memory[1201] = 6'd33;
    assign memory[1202] = 6'd33;
    assign memory[1203] = 6'd33;
    assign memory[1204] = 6'd31;
    assign memory[1205] = 6'd30;
    assign memory[1206] = 6'd29;
    assign memory[1207] = 6'd34;
    assign memory[1208] = 6'd38;
    assign memory[1209] = 6'd37;
    assign memory[1210] = 6'd32;
    assign memory[1211] = 6'd29;
    assign memory[1212] = 6'd29;
    assign memory[1213] = 6'd32;
    assign memory[1214] = 6'd34;
    assign memory[1215] = 6'd33;
    assign memory[1216] = 6'd33;
    assign memory[1217] = 6'd33;
    assign memory[1218] = 6'd33;
    assign memory[1219] = 6'd27;
    assign memory[1220] = 6'd22;
    assign memory[1221] = 6'd24;
    assign memory[1222] = 6'd29;
    assign memory[1223] = 6'd34;
    assign memory[1224] = 6'd33;
    assign memory[1225] = 6'd34;
    assign memory[1226] = 6'd34;
    assign memory[1227] = 6'd34;
    assign memory[1228] = 6'd31;
    assign memory[1229] = 6'd30;
    assign memory[1230] = 6'd30;
    assign memory[1231] = 6'd27;
    assign memory[1232] = 6'd27;
    assign memory[1233] = 6'd27;
    assign memory[1234] = 6'd29;
    assign memory[1235] = 6'd31;
    assign memory[1236] = 6'd31;
    assign memory[1237] = 6'd32;
    assign memory[1238] = 6'd34;
    assign memory[1239] = 6'd34;
    assign memory[1240] = 6'd34;
    assign memory[1241] = 6'd35;
    assign memory[1242] = 6'd34;
    assign memory[1243] = 6'd35;
    assign memory[1244] = 6'd34;
    assign memory[1245] = 6'd33;
    assign memory[1246] = 6'd29;
    assign memory[1247] = 6'd26;
    assign memory[1248] = 6'd27;
    assign memory[1249] = 6'd31;
    assign memory[1250] = 6'd34;
    assign memory[1251] = 6'd33;
    assign memory[1252] = 6'd34;
    assign memory[1253] = 6'd33;
    assign memory[1254] = 6'd33;
    assign memory[1255] = 6'd36;
    assign memory[1256] = 6'd38;
    assign memory[1257] = 6'd37;
    assign memory[1258] = 6'd33;
    assign memory[1259] = 6'd30;
    assign memory[1260] = 6'd30;
    assign memory[1261] = 6'd32;
    assign memory[1262] = 6'd34;
    assign memory[1263] = 6'd33;
    assign memory[1264] = 6'd35;
    assign memory[1265] = 6'd37;
    assign memory[1266] = 6'd37;
    assign memory[1267] = 6'd38;
    assign memory[1268] = 6'd37;
    assign memory[1269] = 6'd37;
    assign memory[1270] = 6'd33;
    assign memory[1271] = 6'd29;
    assign memory[1272] = 6'd31;
    assign memory[1273] = 6'd36;
    assign memory[1274] = 6'd41;
    assign memory[1275] = 6'd39;
    assign memory[1276] = 6'd38;
    assign memory[1277] = 6'd37;
    assign memory[1278] = 6'd37;
    assign memory[1279] = 6'd35;
    assign memory[1280] = 6'd33;
    assign memory[1281] = 6'd34;
    assign memory[1282] = 6'd28;
    assign memory[1283] = 6'd22;
    assign memory[1284] = 6'd23;
    assign memory[1285] = 6'd30;
    assign memory[1286] = 6'd34;
    assign memory[1287] = 6'd34;
    assign memory[1288] = 6'd37;
    assign memory[1289] = 6'd41;
    assign memory[1290] = 6'd40;
    assign memory[1291] = 6'd36;
    assign memory[1292] = 6'd33;
    assign memory[1293] = 6'd34;
    assign memory[1294] = 6'd32;
    assign memory[1295] = 6'd29;
    assign memory[1296] = 6'd30;
    assign memory[1297] = 6'd30;
    assign memory[1298] = 6'd30;
    assign memory[1299] = 6'd30;
    assign memory[1300] = 6'd32;
    assign memory[1301] = 6'd33;
    assign memory[1302] = 6'd33;
    assign memory[1303] = 6'd32;
    assign memory[1304] = 6'd30;
    assign memory[1305] = 6'd30;
    assign memory[1306] = 6'd32;
    assign memory[1307] = 6'd33;
    assign memory[1308] = 6'd33;
    assign memory[1309] = 6'd33;
    assign memory[1310] = 6'd33;
    assign memory[1311] = 6'd34;
    assign memory[1312] = 6'd33;
    assign memory[1313] = 6'd34;
    assign memory[1314] = 6'd33;
    assign memory[1315] = 6'd34;
    assign memory[1316] = 6'd33;
    assign memory[1317] = 6'd33;
    assign memory[1318] = 6'd35;
    assign memory[1319] = 6'd37;
    assign memory[1320] = 6'd37;
    assign memory[1321] = 6'd32;
    assign memory[1322] = 6'd26;
    assign memory[1323] = 6'd26;
    assign memory[1324] = 6'd34;
    assign memory[1325] = 6'd40;
    assign memory[1326] = 6'd40;
    assign memory[1327] = 6'd34;
    assign memory[1328] = 6'd29;
    assign memory[1329] = 6'd30;
    assign memory[1330] = 6'd32;
    assign memory[1331] = 6'd34;
    assign memory[1332] = 6'd34;
    assign memory[1333] = 6'd30;
    assign memory[1334] = 6'd26;
    assign memory[1335] = 6'd26;
    assign memory[1336] = 6'd30;
    assign memory[1337] = 6'd33;
    assign memory[1338] = 6'd34;
    assign memory[1339] = 6'd34;
    assign memory[1340] = 6'd34;
    assign memory[1341] = 6'd34;
    assign memory[1342] = 6'd32;
    assign memory[1343] = 6'd30;
    assign memory[1344] = 6'd30;
    assign memory[1345] = 6'd29;
    assign memory[1346] = 6'd27;
    assign memory[1347] = 6'd26;
    assign memory[1348] = 6'd31;
    assign memory[1349] = 6'd38;
    assign memory[1350] = 6'd38;
    assign memory[1351] = 6'd30;
    assign memory[1352] = 6'd23;
    assign memory[1353] = 6'd23;
    assign memory[1354] = 6'd28;
    assign memory[1355] = 6'd34;
    assign memory[1356] = 6'd35;
    assign memory[1357] = 6'd31;
    assign memory[1358] = 6'd26;
    assign memory[1359] = 6'd26;
    assign memory[1360] = 6'd27;
    assign memory[1361] = 6'd27;
    assign memory[1362] = 6'd27;
    assign memory[1363] = 6'd30;
    assign memory[1364] = 6'd34;
    assign memory[1365] = 6'd34;
    assign memory[1366] = 6'd32;
    assign memory[1367] = 6'd30;
    assign memory[1368] = 6'd29;
    assign memory[1369] = 6'd28;
    assign memory[1370] = 6'd27;
    assign memory[1371] = 6'd27;
    assign memory[1372] = 6'd29;
    assign memory[1373] = 6'd30;
    assign memory[1374] = 6'd30;
    assign memory[1375] = 6'd30;
    assign memory[1376] = 6'd31;
    assign memory[1377] = 6'd30;
    assign memory[1378] = 6'd30;
    assign memory[1379] = 6'd30;
    assign memory[1380] = 6'd29;
    assign memory[1381] = 6'd33;
    assign memory[1382] = 6'd37;
    assign memory[1383] = 6'd37;
    assign memory[1384] = 6'd33;
    assign memory[1385] = 6'd27;
    assign memory[1386] = 6'd27;
    assign memory[1387] = 6'd28;
    assign memory[1388] = 6'd31;
    assign memory[1389] = 6'd30;
    assign memory[1390] = 6'd30;
    assign memory[1391] = 6'd31;
    assign memory[1392] = 6'd30;
    assign memory[1393] = 6'd32;
    assign memory[1394] = 6'd33;
    assign memory[1395] = 6'd34;
    assign memory[1396] = 6'd30;
    assign memory[1397] = 6'd23;
    assign memory[1398] = 6'd23;
    assign memory[1399] = 6'd30;
    assign memory[1400] = 6'd37;
    assign memory[1401] = 6'd37;
    assign memory[1402] = 6'd32;
    assign memory[1403] = 6'd26;
    assign memory[1404] = 6'd27;
    assign memory[1405] = 6'd30;
    assign memory[1406] = 6'd31;
    assign memory[1407] = 6'd30;
    assign memory[1408] = 6'd31;
    assign memory[1409] = 6'd34;
    assign memory[1410] = 6'd33;
    assign memory[1411] = 6'd35;
    assign memory[1412] = 6'd37;
    assign memory[1413] = 6'd38;
    assign memory[1414] = 6'd34;
    assign memory[1415] = 6'd30;
    assign memory[1416] = 6'd29;
    assign memory[1417] = 6'd33;
    assign memory[1418] = 6'd37;
    assign memory[1419] = 6'd37;
    assign memory[1420] = 6'd36;
    assign memory[1421] = 6'd37;
    assign memory[1422] = 6'd37;
    assign memory[1423] = 6'd37;
    assign memory[1424] = 6'd36;
    assign memory[1425] = 6'd36;
    assign memory[1426] = 6'd37;
    assign memory[1427] = 6'd36;
    assign memory[1428] = 6'd36;
    assign memory[1429] = 6'd35;
    assign memory[1430] = 6'd32;
    assign memory[1431] = 6'd32;
    assign memory[1432] = 6'd34;
    assign memory[1433] = 6'd36;
    assign memory[1434] = 6'd37;
    assign memory[1435] = 6'd35;
    assign memory[1436] = 6'd34;
    assign memory[1437] = 6'd34;
    assign memory[1438] = 6'd32;
    assign memory[1439] = 6'd30;
    assign memory[1440] = 6'd29;
    assign memory[1441] = 6'd31;
    assign memory[1442] = 6'd32;
    assign memory[1443] = 6'd33;
    assign memory[1444] = 6'd35;
    assign memory[1445] = 6'd36;
    assign memory[1446] = 6'd37;
    assign memory[1447] = 6'd33;
    assign memory[1448] = 6'd30;
    assign memory[1449] = 6'd29;
    assign memory[1450] = 6'd31;
    assign memory[1451] = 6'd33;
    assign memory[1452] = 6'd34;
    assign memory[1453] = 6'd33;
    assign memory[1454] = 6'd34;
    assign memory[1455] = 6'd34;
    assign memory[1456] = 6'd34;
    assign memory[1457] = 6'd34;
    assign memory[1458] = 6'd33;
    assign memory[1459] = 6'd33;
    assign memory[1460] = 6'd33;
    assign memory[1461] = 6'd34;
    assign memory[1462] = 6'd32;
    assign memory[1463] = 6'd30;
    assign memory[1464] = 6'd30;
    assign memory[1465] = 6'd29;
    assign memory[1466] = 6'd27;
    assign memory[1467] = 6'd26;
    assign memory[1468] = 6'd31;
    assign memory[1469] = 6'd37;
    assign memory[1470] = 6'd37;
    assign memory[1471] = 6'd34;
    assign memory[1472] = 6'd30;
    assign memory[1473] = 6'd29;
    assign memory[1474] = 6'd33;
    assign memory[1475] = 6'd37;
    assign memory[1476] = 6'd38;
    assign memory[1477] = 6'd37;
    assign memory[1478] = 6'd37;
    assign memory[1479] = 6'd37;
    assign memory[1480] = 6'd37;
    assign memory[1481] = 6'd36;
    assign memory[1482] = 6'd37;
    assign memory[1483] = 6'd34;
    assign memory[1484] = 6'd30;
    assign memory[1485] = 6'd30;
    assign memory[1486] = 6'd33;
    assign memory[1487] = 6'd37;
    assign memory[1488] = 6'd38;
    assign memory[1489] = 6'd34;
    assign memory[1490] = 6'd30;
    assign memory[1491] = 6'd30;
    assign memory[1492] = 6'd33;
    assign memory[1493] = 6'd37;
    assign memory[1494] = 6'd37;
    assign memory[1495] = 6'd35;
    assign memory[1496] = 6'd34;
    assign memory[1497] = 6'd33;
    assign memory[1498] = 6'd33;
    assign memory[1499] = 6'd33;
    assign memory[1500] = 6'd33;
    assign memory[1501] = 6'd32;
    assign memory[1502] = 6'd30;
    assign memory[1503] = 6'd30;
    assign memory[1504] = 6'd30;
    assign memory[1505] = 6'd31;
    assign memory[1506] = 6'd31;
    assign memory[1507] = 6'd31;
    assign memory[1508] = 6'd30;
    assign memory[1509] = 6'd30;
    assign memory[1510] = 6'd31;
    assign memory[1511] = 6'd34;
    assign memory[1512] = 6'd33;
    assign memory[1513] = 6'd33;
    assign memory[1514] = 6'd32;
    assign memory[1515] = 6'd33;
    assign memory[1516] = 6'd32;
    assign memory[1517] = 6'd30;
    assign memory[1518] = 6'd31;
    assign memory[1519] = 6'd31;
    assign memory[1520] = 6'd31;
    assign memory[1521] = 6'd30;
    assign memory[1522] = 6'd31;
    assign memory[1523] = 6'd33;
    assign memory[1524] = 6'd33;
    assign memory[1525] = 6'd33;
    assign memory[1526] = 6'd33;
    assign memory[1527] = 6'd33;
    assign memory[1528] = 6'd29;
    assign memory[1529] = 6'd20;
    assign memory[1530] = 6'd18;
    assign memory[1531] = 6'd25;
    assign memory[1532] = 6'd33;
    assign memory[1533] = 6'd35;
    assign memory[1534] = 6'd31;
    assign memory[1535] = 6'd26;
    assign memory[1536] = 6'd26;
    assign memory[1537] = 6'd28;
    assign memory[1538] = 6'd30;
    assign memory[1539] = 6'd31;
    assign memory[1540] = 6'd28;
    assign memory[1541] = 6'd27;
    assign memory[1542] = 6'd26;
    assign memory[1543] = 6'd28;
    assign memory[1544] = 6'd29;
    assign memory[1545] = 6'd30;
    assign memory[1546] = 6'd30;
    assign memory[1547] = 6'd30;
    assign memory[1548] = 6'd32;
    assign memory[1549] = 6'd30;
    assign memory[1550] = 6'd27;
    assign memory[1551] = 6'd27;
    assign memory[1552] = 6'd27;
    assign memory[1553] = 6'd27;
    assign memory[1554] = 6'd26;
    assign memory[1555] = 6'd29;
    assign memory[1556] = 6'd34;
    assign memory[1557] = 6'd34;
    assign memory[1558] = 6'd33;
    assign memory[1559] = 6'd29;
    assign memory[1560] = 6'd30;
    assign memory[1561] = 6'd29;
    assign memory[1562] = 6'd27;
    assign memory[1563] = 6'd26;
    assign memory[1564] = 6'd28;
    assign memory[1565] = 6'd33;
    assign memory[1566] = 6'd34;
    assign memory[1567] = 6'd33;
    assign memory[1568] = 6'd30;
    assign memory[1569] = 6'd30;
    assign memory[1570] = 6'd31;
    assign memory[1571] = 6'd30;
    assign memory[1572] = 6'd30;
    assign memory[1573] = 6'd30;
    assign memory[1574] = 6'd30;
    assign memory[1575] = 6'd29;
    assign memory[1576] = 6'd30;
    assign memory[1577] = 6'd30;
    assign memory[1578] = 6'd30;
    assign memory[1579] = 6'd29;
    assign memory[1580] = 6'd30;
    assign memory[1581] = 6'd30;
    assign memory[1582] = 6'd31;
    assign memory[1583] = 6'd36;
    assign memory[1584] = 6'd37;
    assign memory[1585] = 6'd34;
    assign memory[1586] = 6'd27;
    assign memory[1587] = 6'd26;
    assign memory[1588] = 6'd30;
    assign memory[1589] = 6'd37;
    assign memory[1590] = 6'd38;
    assign memory[1591] = 6'd33;
    assign memory[1592] = 6'd27;
    assign memory[1593] = 6'd25;
    assign memory[1594] = 6'd28;
    assign memory[1595] = 6'd32;
    assign memory[1596] = 6'd34;
    assign memory[1597] = 6'd32;
    assign memory[1598] = 6'd30;
    assign memory[1599] = 6'd30;
    assign memory[1600] = 6'd30;
    assign memory[1601] = 6'd30;
    assign memory[1602] = 6'd30;
    assign memory[1603] = 6'd31;
    assign memory[1604] = 6'd34;
    assign memory[1605] = 6'd34;
    assign memory[1606] = 6'd34;
    assign memory[1607] = 6'd36;
    assign memory[1608] = 6'd36;
    assign memory[1609] = 6'd36;
    assign memory[1610] = 6'd33;
    assign memory[1611] = 6'd33;
    assign memory[1612] = 6'd32;
    assign memory[1613] = 6'd30;
    assign memory[1614] = 6'd30;
    assign memory[1615] = 6'd31;
    assign memory[1616] = 6'd30;
    assign memory[1617] = 6'd30;
    assign memory[1618] = 6'd30;
    assign memory[1619] = 6'd30;
    assign memory[1620] = 6'd30;
    assign memory[1621] = 6'd30;
    assign memory[1622] = 6'd30;
    assign memory[1623] = 6'd29;
    assign memory[1624] = 6'd30;
    assign memory[1625] = 6'd33;
    assign memory[1626] = 6'd34;
    assign memory[1627] = 6'd33;
    assign memory[1628] = 6'd34;
    assign memory[1629] = 6'd33;
    assign memory[1630] = 6'd33;
    assign memory[1631] = 6'd30;
    assign memory[1632] = 6'd29;
    assign memory[1633] = 6'd32;
    assign memory[1634] = 6'd36;
    assign memory[1635] = 6'd37;
    assign memory[1636] = 6'd35;
    assign memory[1637] = 6'd34;
    assign memory[1638] = 6'd33;
    assign memory[1639] = 6'd34;
    assign memory[1640] = 6'd34;
    assign memory[1641] = 6'd34;
    assign memory[1642] = 6'd34;
    assign memory[1643] = 6'd34;
    assign memory[1644] = 6'd34;
    assign memory[1645] = 6'd33;
    assign memory[1646] = 6'd33;
    assign memory[1647] = 6'd33;
    assign memory[1648] = 6'd33;
    assign memory[1649] = 6'd33;
    assign memory[1650] = 6'd34;
    assign memory[1651] = 6'd33;
    assign memory[1652] = 6'd30;
    assign memory[1653] = 6'd29;
    assign memory[1654] = 6'd31;
    assign memory[1655] = 6'd33;
    assign memory[1656] = 6'd34;
    assign memory[1657] = 6'd33;
    assign memory[1658] = 6'd31;
    assign memory[1659] = 6'd30;
    assign memory[1660] = 6'd30;
    assign memory[1661] = 6'd33;
    assign memory[1662] = 6'd34;
    assign memory[1663] = 6'd33;
    assign memory[1664] = 6'd31;
    assign memory[1665] = 6'd30;
    assign memory[1666] = 6'd30;
    assign memory[1667] = 6'd30;
    assign memory[1668] = 6'd30;
    assign memory[1669] = 6'd30;
    assign memory[1670] = 6'd30;
    assign memory[1671] = 6'd30;
    assign memory[1672] = 6'd31;
    assign memory[1673] = 6'd33;
    assign memory[1674] = 6'd33;
    assign memory[1675] = 6'd33;
    assign memory[1676] = 6'd34;
    assign memory[1677] = 6'd34;
    assign memory[1678] = 6'd33;
    assign memory[1679] = 6'd31;
    assign memory[1680] = 6'd30;
    assign memory[1681] = 6'd30;
    assign memory[1682] = 6'd31;
    assign memory[1683] = 6'd31;
    assign memory[1684] = 6'd31;
    assign memory[1685] = 6'd30;
    assign memory[1686] = 6'd30;
    assign memory[1687] = 6'd30;
    assign memory[1688] = 6'd30;
    assign memory[1689] = 6'd30;
    assign memory[1690] = 6'd32;
    assign memory[1691] = 6'd34;
    assign memory[1692] = 6'd35;
    assign memory[1693] = 6'd33;
    assign memory[1694] = 6'd30;
    assign memory[1695] = 6'd30;
    assign memory[1696] = 6'd30;
    assign memory[1697] = 6'd29;
    assign memory[1698] = 6'd30;
    assign memory[1699] = 6'd31;
    assign memory[1700] = 6'd33;
    assign memory[1701] = 6'd33;
    assign memory[1702] = 6'd33;
    assign memory[1703] = 6'd30;
    assign memory[1704] = 6'd30;
    assign memory[1705] = 6'd30;
    assign memory[1706] = 6'd27;
    assign memory[1707] = 6'd26;
    assign memory[1708] = 6'd27;
    assign memory[1709] = 6'd30;
    assign memory[1710] = 6'd30;
    assign memory[1711] = 6'd31;
    assign memory[1712] = 6'd30;
    assign memory[1713] = 6'd30;
    assign memory[1714] = 6'd31;
    assign memory[1715] = 6'd33;
    assign memory[1716] = 6'd34;
    assign memory[1717] = 6'd33;
    assign memory[1718] = 6'd33;
    assign memory[1719] = 6'd33;
    assign memory[1720] = 6'd32;
    assign memory[1721] = 6'd30;
    assign memory[1722] = 6'd30;
    assign memory[1723] = 6'd30;
    assign memory[1724] = 6'd30;
    assign memory[1725] = 6'd30;
    assign memory[1726] = 6'd30;
    assign memory[1727] = 6'd29;
    assign memory[1728] = 6'd29;
    assign memory[1729] = 6'd29;
    assign memory[1730] = 6'd30;
    assign memory[1731] = 6'd29;
    assign memory[1732] = 6'd31;
    assign memory[1733] = 6'd33;
    assign memory[1734] = 6'd34;
    assign memory[1735] = 6'd32;
    assign memory[1736] = 6'd30;
    assign memory[1737] = 6'd29;
    assign memory[1738] = 6'd30;
    assign memory[1739] = 6'd30;
    assign memory[1740] = 6'd30;
    assign memory[1741] = 6'd30;
    assign memory[1742] = 6'd32;
    assign memory[1743] = 6'd33;
    assign memory[1744] = 6'd33;
    assign memory[1745] = 6'd33;
    assign memory[1746] = 6'd34;
    assign memory[1747] = 6'd33;
    assign memory[1748] = 6'd31;
    assign memory[1749] = 6'd30;
    assign memory[1750] = 6'd31;
    assign memory[1751] = 6'd33;
    assign memory[1752] = 6'd33;
    assign memory[1753] = 6'd33;
    assign memory[1754] = 6'd33;
    assign memory[1755] = 6'd33;
    assign memory[1756] = 6'd33;
    assign memory[1757] = 6'd30;
    assign memory[1758] = 6'd29;
    assign memory[1759] = 6'd31;
    assign memory[1760] = 6'd36;
    assign memory[1761] = 6'd38;
    assign memory[1762] = 6'd35;
    assign memory[1763] = 6'd31;
    assign memory[1764] = 6'd29;
    assign memory[1765] = 6'd31;
    assign memory[1766] = 6'd33;
    assign memory[1767] = 6'd34;
    assign memory[1768] = 6'd33;
    assign memory[1769] = 6'd31;
    assign memory[1770] = 6'd30;
    assign memory[1771] = 6'd31;
    assign memory[1772] = 6'd35;
    assign memory[1773] = 6'd37;
    assign memory[1774] = 6'd36;
    assign memory[1775] = 6'd30;
    assign memory[1776] = 6'd30;
    assign memory[1777] = 6'd29;
    assign memory[1778] = 6'd27;
    assign memory[1779] = 6'd27;
    assign memory[1780] = 6'd28;
    assign memory[1781] = 6'd30;
    assign memory[1782] = 6'd30;
    assign memory[1783] = 6'd30;
    assign memory[1784] = 6'd33;
    assign memory[1785] = 6'd33;
    assign memory[1786] = 6'd33;
    assign memory[1787] = 6'd31;
    assign memory[1788] = 6'd30;
    assign memory[1789] = 6'd31;
    assign memory[1790] = 6'd33;
    assign memory[1791] = 6'd35;
    assign memory[1792] = 6'd33;
    assign memory[1793] = 6'd28;
    assign memory[1794] = 6'd25;
    assign memory[1795] = 6'd27;
    assign memory[1796] = 6'd32;
    assign memory[1797] = 6'd34;
    assign memory[1798] = 6'd33;
    assign memory[1799] = 6'd30;
    assign memory[1800] = 6'd29;
    assign memory[1801] = 6'd30;
    assign memory[1802] = 6'd33;
    assign memory[1803] = 6'd34;
    assign memory[1804] = 6'd33;
    assign memory[1805] = 6'd31;
    assign memory[1806] = 6'd30;
    assign memory[1807] = 6'd31;
    assign memory[1808] = 6'd30;
    assign memory[1809] = 6'd29;
    assign memory[1810] = 6'd31;
    assign memory[1811] = 6'd33;
    assign memory[1812] = 6'd34;
    assign memory[1813] = 6'd33;
    assign memory[1814] = 6'd31;
    assign memory[1815] = 6'd30;
    assign memory[1816] = 6'd30;
    assign memory[1817] = 6'd30;
    assign memory[1818] = 6'd31;
    assign memory[1819] = 6'd30;
    assign memory[1820] = 6'd31;
    assign memory[1821] = 6'd30;
    assign memory[1822] = 6'd30;
    assign memory[1823] = 6'd32;
    assign memory[1824] = 6'd34;
    assign memory[1825] = 6'd34;
    assign memory[1826] = 6'd34;
    assign memory[1827] = 6'd33;
    assign memory[1828] = 6'd33;
    assign memory[1829] = 6'd30;
    assign memory[1830] = 6'd29;
    assign memory[1831] = 6'd30;
    assign memory[1832] = 6'd29;
    assign memory[1833] = 6'd30;
    assign memory[1834] = 6'd31;
    assign memory[1835] = 6'd32;
    assign memory[1836] = 6'd34;
    assign memory[1837] = 6'd33;
    assign memory[1838] = 6'd31;
    assign memory[1839] = 6'd30;
    assign memory[1840] = 6'd30;
    assign memory[1841] = 6'd32;
    assign memory[1842] = 6'd34;
    assign memory[1843] = 6'd33;
    assign memory[1844] = 6'd31;
    assign memory[1845] = 6'd30;
    assign memory[1846] = 6'd31;
    assign memory[1847] = 6'd33;
    assign memory[1848] = 6'd33;
    assign memory[1849] = 6'd33;
    assign memory[1850] = 6'd33;
    assign memory[1851] = 6'd34;
    assign memory[1852] = 6'd33;
    assign memory[1853] = 6'd31;
    assign memory[1854] = 6'd29;
    assign memory[1855] = 6'd30;
    assign memory[1856] = 6'd33;
    assign memory[1857] = 6'd33;
    assign memory[1858] = 6'd33;
    assign memory[1859] = 6'd30;
    assign memory[1860] = 6'd30;
    assign memory[1861] = 6'd30;
    assign memory[1862] = 6'd31;
    assign memory[1863] = 6'd30;
    assign memory[1864] = 6'd30;
    assign memory[1865] = 6'd32;
    assign memory[1866] = 6'd33;
    assign memory[1867] = 6'd33;
    assign memory[1868] = 6'd30;
    assign memory[1869] = 6'd30;
    assign memory[1870] = 6'd29;
    assign memory[1871] = 6'd27;
    assign memory[1872] = 6'd27;
    assign memory[1873] = 6'd27;
    assign memory[1874] = 6'd30;
    assign memory[1875] = 6'd31;
    assign memory[1876] = 6'd30;
    assign memory[1877] = 6'd32;
    assign memory[1878] = 6'd34;
    assign memory[1879] = 6'd33;
    assign memory[1880] = 6'd31;
    assign memory[1881] = 6'd29;
    assign memory[1882] = 6'd30;
    assign memory[1883] = 6'd29;
    assign memory[1884] = 6'd30;
    assign memory[1885] = 6'd30;
    assign memory[1886] = 6'd30;
    assign memory[1887] = 6'd30;
    assign memory[1888] = 6'd30;
    assign memory[1889] = 6'd33;
    assign memory[1890] = 6'd34;
    assign memory[1891] = 6'd33;
    assign memory[1892] = 6'd32;
    assign memory[1893] = 6'd30;
    assign memory[1894] = 6'd30;
    assign memory[1895] = 6'd29;
    assign memory[1896] = 6'd29;
    assign memory[1897] = 6'd29;
    assign memory[1898] = 6'd29;
    assign memory[1899] = 6'd29;
    assign memory[1900] = 6'd29;
    assign memory[1901] = 6'd33;
    assign memory[1902] = 6'd34;
    assign memory[1903] = 6'd34;
    assign memory[1904] = 6'd34;
    assign memory[1905] = 6'd34;
    assign memory[1906] = 6'd33;
    assign memory[1907] = 6'd31;
    assign memory[1908] = 6'd30;
    assign memory[1909] = 6'd31;
    assign memory[1910] = 6'd33;
    assign memory[1911] = 6'd34;
    assign memory[1912] = 6'd33;
    assign memory[1913] = 6'd31;
    assign memory[1914] = 6'd30;
    assign memory[1915] = 6'd30;
    assign memory[1916] = 6'd30;
    assign memory[1917] = 6'd30;
    assign memory[1918] = 6'd31;
    assign memory[1919] = 6'd33;
    assign memory[1920] = 6'd34;
    assign memory[1921] = 6'd34;
    assign memory[1922] = 6'd34;
    assign memory[1923] = 6'd34;
    assign memory[1924] = 6'd33;
    assign memory[1925] = 6'd31;
    assign memory[1926] = 6'd29;
    assign memory[1927] = 6'd30;
    assign memory[1928] = 6'd33;
    assign memory[1929] = 6'd34;
    assign memory[1930] = 6'd33;
    assign memory[1931] = 6'd31;
    assign memory[1932] = 6'd30;
    assign memory[1933] = 6'd31;
    assign memory[1934] = 6'd33;
    assign memory[1935] = 6'd34;
    assign memory[1936] = 6'd33;
    assign memory[1937] = 6'd31;
    assign memory[1938] = 6'd29;
    assign memory[1939] = 6'd30;
    assign memory[1940] = 6'd32;
    assign memory[1941] = 6'd34;
    assign memory[1942] = 6'd33;
    assign memory[1943] = 6'd32;
    assign memory[1944] = 6'd30;
    assign memory[1945] = 6'd30;
    assign memory[1946] = 6'd30;
    assign memory[1947] = 6'd30;
    assign memory[1948] = 6'd30;
    assign memory[1949] = 6'd28;
    assign memory[1950] = 6'd26;
    assign memory[1951] = 6'd27;
    assign memory[1952] = 6'd31;
    assign memory[1953] = 6'd34;
    assign memory[1954] = 6'd34;
    assign memory[1955] = 6'd34;
    assign memory[1956] = 6'd34;
    assign memory[1957] = 6'd33;
    assign memory[1958] = 6'd31;
    assign memory[1959] = 6'd30;
    assign memory[1960] = 6'd31;
    assign memory[1961] = 6'd30;
    assign memory[1962] = 6'd30;
    assign memory[1963] = 6'd30;
    assign memory[1964] = 6'd31;
    assign memory[1965] = 6'd30;
    assign memory[1966] = 6'd31;
    assign memory[1967] = 6'd33;
    assign memory[1968] = 6'd34;
    assign memory[1969] = 6'd34;
    assign memory[1970] = 6'd31;
    assign memory[1971] = 6'd30;
    assign memory[1972] = 6'd30;
    assign memory[1973] = 6'd33;
    assign memory[1974] = 6'd34;
    assign memory[1975] = 6'd33;
    assign memory[1976] = 6'd31;
    assign memory[1977] = 6'd29;
    assign memory[1978] = 6'd30;
    assign memory[1979] = 6'd30;
    assign memory[1980] = 6'd30;
    assign memory[1981] = 6'd30;
    assign memory[1982] = 6'd30;
    assign memory[1983] = 6'd30;
    assign memory[1984] = 6'd30;
    assign memory[1985] = 6'd30;
    assign memory[1986] = 6'd30;
    assign memory[1987] = 6'd30;
    assign memory[1988] = 6'd28;
    assign memory[1989] = 6'd25;
    assign memory[1990] = 6'd27;
    assign memory[1991] = 6'd30;
    assign memory[1992] = 6'd34;
    assign memory[1993] = 6'd33;
    assign memory[1994] = 6'd26;
    assign memory[1995] = 6'd22;
    assign memory[1996] = 6'd23;
    assign memory[1997] = 6'd28;
    assign memory[1998] = 6'd31;
    assign memory[1999] = 6'd29;
    assign memory[2000] = 6'd27;
    assign memory[2001] = 6'd25;
    assign memory[2002] = 6'd27;
    assign memory[2003] = 6'd31;
    assign memory[2004] = 6'd34;
    assign memory[2005] = 6'd33;
    assign memory[2006] = 6'd33;
    assign memory[2007] = 6'd34;
    assign memory[2008] = 6'd34;
    assign memory[2009] = 6'd30;
    assign memory[2010] = 6'd26;
    assign memory[2011] = 6'd27;
    assign memory[2012] = 6'd31;
    assign memory[2013] = 6'd35;
    assign memory[2014] = 6'd33;
    assign memory[2015] = 6'd30;
    assign memory[2016] = 6'd26;
    assign memory[2017] = 6'd27;
    assign memory[2018] = 6'd30;
    assign memory[2019] = 6'd34;
    assign memory[2020] = 6'd33;
    assign memory[2021] = 6'd31;
    assign memory[2022] = 6'd30;
    assign memory[2023] = 6'd31;
    assign memory[2024] = 6'd33;
    assign memory[2025] = 6'd34;
    assign memory[2026] = 6'd34;
    assign memory[2027] = 6'd33;
    assign memory[2028] = 6'd34;
    assign memory[2029] = 6'd33;
    assign memory[2030] = 6'd33;
    assign memory[2031] = 6'd33;
    assign memory[2032] = 6'd33;
    assign memory[2033] = 6'd34;
    assign memory[2034] = 6'd34;
    assign memory[2035] = 6'd34;
    assign memory[2036] = 6'd34;
    assign memory[2037] = 6'd34;
    assign memory[2038] = 6'd33;
    assign memory[2039] = 6'd34;
    assign memory[2040] = 6'd32;
    assign memory[2041] = 6'd34;
    assign memory[2042] = 6'd35;
    assign memory[2043] = 6'd37;
    assign memory[2044] = 6'd36;
    assign memory[2045] = 6'd32;
    assign memory[2046] = 6'd29;
    assign memory[2047] = 6'd30;
    assign memory[2048] = 6'd32;
    assign memory[2049] = 6'd34;
    assign memory[2050] = 6'd33;
    assign memory[2051] = 6'd31;
    assign memory[2052] = 6'd30;
    assign memory[2053] = 6'd30;
    assign memory[2054] = 6'd32;
    assign memory[2055] = 6'd33;
    assign memory[2056] = 6'd33;
    assign memory[2057] = 6'd33;
    assign memory[2058] = 6'd33;
    assign memory[2059] = 6'd32;
    assign memory[2060] = 6'd33;
    assign memory[2061] = 6'd33;
    assign memory[2062] = 6'd34;
    assign memory[2063] = 6'd33;
    assign memory[2064] = 6'd33;
    assign memory[2065] = 6'd34;
    assign memory[2066] = 6'd32;
    assign memory[2067] = 6'd30;
    assign memory[2068] = 6'd30;
    assign memory[2069] = 6'd32;
    assign memory[2070] = 6'd34;
    assign memory[2071] = 6'd34;
    assign memory[2072] = 6'd30;
    assign memory[2073] = 6'd26;
    assign memory[2074] = 6'd26;
    assign memory[2075] = 6'd31;
    assign memory[2076] = 6'd34;
    assign memory[2077] = 6'd33;
    assign memory[2078] = 6'd31;
    assign memory[2079] = 6'd29;
    assign memory[2080] = 6'd30;
    assign memory[2081] = 6'd32;
    assign memory[2082] = 6'd34;
    assign memory[2083] = 6'd34;
    assign memory[2084] = 6'd34;
    assign memory[2085] = 6'd34;
    assign memory[2086] = 6'd34;
    assign memory[2087] = 6'd34;
    assign memory[2088] = 6'd34;
    assign memory[2089] = 6'd34;
    assign memory[2090] = 6'd31;
    assign memory[2091] = 6'd31;
    assign memory[2092] = 6'd30;
    assign memory[2093] = 6'd31;
    assign memory[2094] = 6'd30;
    assign memory[2095] = 6'd30;
    assign memory[2096] = 6'd30;
    assign memory[2097] = 6'd30;
    assign memory[2098] = 6'd31;
    assign memory[2099] = 6'd31;
    assign memory[2100] = 6'd30;
    assign memory[2101] = 6'd31;
    assign memory[2102] = 6'd33;
    assign memory[2103] = 6'd34;
    assign memory[2104] = 6'd34;
    assign memory[2105] = 6'd32;
    assign memory[2106] = 6'd31;
    assign memory[2107] = 6'd31;
    assign memory[2108] = 6'd29;
    assign memory[2109] = 6'd27;
    assign memory[2110] = 6'd26;
    assign memory[2111] = 6'd29;
    assign memory[2112] = 6'd30;
    assign memory[2113] = 6'd30;
    assign memory[2114] = 6'd31;
    assign memory[2115] = 6'd31;
    assign memory[2116] = 6'd31;
    assign memory[2117] = 6'd30;
    assign memory[2118] = 6'd30;
    assign memory[2119] = 6'd30;
    assign memory[2120] = 6'd30;
    assign memory[2121] = 6'd30;
    assign memory[2122] = 6'd30;
    assign memory[2123] = 6'd31;
    assign memory[2124] = 6'd30;
    assign memory[2125] = 6'd30;
    assign memory[2126] = 6'd30;
    assign memory[2127] = 6'd31;
    assign memory[2128] = 6'd30;
    assign memory[2129] = 6'd30;
    assign memory[2130] = 6'd31;
    assign memory[2131] = 6'd30;
    assign memory[2132] = 6'd31;
    assign memory[2133] = 6'd31;
    assign memory[2134] = 6'd31;
    assign memory[2135] = 6'd31;
    assign memory[2136] = 6'd31;
    assign memory[2137] = 6'd30;
    assign memory[2138] = 6'd31;
    assign memory[2139] = 6'd34;
    assign memory[2140] = 6'd34;
    assign memory[2141] = 6'd32;
    assign memory[2142] = 6'd30;
    assign memory[2143] = 6'd30;
    assign memory[2144] = 6'd32;
    assign memory[2145] = 6'd33;
    assign memory[2146] = 6'd33;
    assign memory[2147] = 6'd32;
    assign memory[2148] = 6'd30;
    assign memory[2149] = 6'd30;
    assign memory[2150] = 6'd32;
    assign memory[2151] = 6'd33;
    assign memory[2152] = 6'd33;
    assign memory[2153] = 6'd34;
    assign memory[2154] = 6'd34;
    assign memory[2155] = 6'd34;
    assign memory[2156] = 6'd32;
    assign memory[2157] = 6'd30;
    assign memory[2158] = 6'd29;
    assign memory[2159] = 6'd32;
    assign memory[2160] = 6'd34;
    assign memory[2161] = 6'd34;
    assign memory[2162] = 6'd32;
    assign memory[2163] = 6'd30;
    assign memory[2164] = 6'd30;
    assign memory[2165] = 6'd31;
    assign memory[2166] = 6'd30;
    assign memory[2167] = 6'd30;
    assign memory[2168] = 6'd32;
    assign memory[2169] = 6'd34;
    assign memory[2170] = 6'd33;
    assign memory[2171] = 6'd32;
    assign memory[2172] = 6'd30;
    assign memory[2173] = 6'd30;
    assign memory[2174] = 6'd30;
    assign memory[2175] = 6'd30;
    assign memory[2176] = 6'd30;
    assign memory[2177] = 6'd30;
    assign memory[2178] = 6'd30;
    assign memory[2179] = 6'd30;
    assign memory[2180] = 6'd32;
    assign memory[2181] = 6'd34;
    assign memory[2182] = 6'd34;
    assign memory[2183] = 6'd30;
    assign memory[2184] = 6'd26;
    assign memory[2185] = 6'd27;
    assign memory[2186] = 6'd29;
    assign memory[2187] = 6'd31;
    assign memory[2188] = 6'd30;
    assign memory[2189] = 6'd31;
    assign memory[2190] = 6'd30;
    assign memory[2191] = 6'd30;
    assign memory[2192] = 6'd32;
    assign memory[2193] = 6'd34;
    assign memory[2194] = 6'd34;
    assign memory[2195] = 6'd32;
    assign memory[2196] = 6'd30;
    assign memory[2197] = 6'd30;
    assign memory[2198] = 6'd32;
    assign memory[2199] = 6'd33;
    assign memory[2200] = 6'd33;
    assign memory[2201] = 6'd32;
    assign memory[2202] = 6'd29;
    assign memory[2203] = 6'd29;
    assign memory[2204] = 6'd30;
    assign memory[2205] = 6'd30;
    assign memory[2206] = 6'd30;
    assign memory[2207] = 6'd32;
    assign memory[2208] = 6'd33;
    assign memory[2209] = 6'd33;
    assign memory[2210] = 6'd33;
    assign memory[2211] = 6'd34;
    assign memory[2212] = 6'd34;
    assign memory[2213] = 6'd33;
    assign memory[2214] = 6'd33;
    assign memory[2215] = 6'd34;
    assign memory[2216] = 6'd34;
    assign memory[2217] = 6'd33;
    assign memory[2218] = 6'd33;
    assign memory[2219] = 6'd33;
    assign memory[2220] = 6'd33;
    assign memory[2221] = 6'd34;
    assign memory[2222] = 6'd33;
    assign memory[2223] = 6'd33;
    assign memory[2224] = 6'd33;
    assign memory[2225] = 6'd33;
    assign memory[2226] = 6'd33;
    assign memory[2227] = 6'd33;
    assign memory[2228] = 6'd32;
    assign memory[2229] = 6'd30;
    assign memory[2230] = 6'd30;
    assign memory[2231] = 6'd32;
    assign memory[2232] = 6'd34;
    assign memory[2233] = 6'd34;
    assign memory[2234] = 6'd31;
    assign memory[2235] = 6'd30;
    assign memory[2236] = 6'd30;
    assign memory[2237] = 6'd32;
    assign memory[2238] = 6'd34;
    assign memory[2239] = 6'd34;
    assign memory[2240] = 6'd32;
    assign memory[2241] = 6'd30;
    assign memory[2242] = 6'd30;
    assign memory[2243] = 6'd31;
    assign memory[2244] = 6'd31;
    assign memory[2245] = 6'd30;
    assign memory[2246] = 6'd32;
    assign memory[2247] = 6'd34;
    assign memory[2248] = 6'd34;
    assign memory[2249] = 6'd34;
    assign memory[2250] = 6'd33;
    assign memory[2251] = 6'd33;
    assign memory[2252] = 6'd32;
    assign memory[2253] = 6'd30;
    assign memory[2254] = 6'd29;
    assign memory[2255] = 6'd32;
    assign memory[2256] = 6'd34;
    assign memory[2257] = 6'd34;
    assign memory[2258] = 6'd33;
    assign memory[2259] = 6'd33;
    assign memory[2260] = 6'd33;
    assign memory[2261] = 6'd32;
    assign memory[2262] = 6'd30;
    assign memory[2263] = 6'd30;
    assign memory[2264] = 6'd32;
    assign memory[2265] = 6'd34;
    assign memory[2266] = 6'd34;
    assign memory[2267] = 6'd34;
    assign memory[2268] = 6'd33;
    assign memory[2269] = 6'd34;
    assign memory[2270] = 6'd32;
    assign memory[2271] = 6'd30;
    assign memory[2272] = 6'd30;
    assign memory[2273] = 6'd30;
    assign memory[2274] = 6'd31;
    assign memory[2275] = 6'd30;
    assign memory[2276] = 6'd31;
    assign memory[2277] = 6'd34;
    assign memory[2278] = 6'd33;
    assign memory[2279] = 6'd32;
    assign memory[2280] = 6'd31;
    assign memory[2281] = 6'd31;
    assign memory[2282] = 6'd30;
    assign memory[2283] = 6'd30;
    assign memory[2284] = 6'd31;
    assign memory[2285] = 6'd31;
    assign memory[2286] = 6'd31;
    assign memory[2287] = 6'd30;
    assign memory[2288] = 6'd31;
    assign memory[2289] = 6'd34;
    assign memory[2290] = 6'd34;
    assign memory[2291] = 6'd33;
    assign memory[2292] = 6'd31;
    assign memory[2293] = 6'd30;
    assign memory[2294] = 6'd30;
    assign memory[2295] = 6'd30;
    assign memory[2296] = 6'd30;
    assign memory[2297] = 6'd30;
    assign memory[2298] = 6'd30;
    assign memory[2299] = 6'd30;
    assign memory[2300] = 6'd31;
    assign memory[2301] = 6'd31;
    assign memory[2302] = 6'd30;
    assign memory[2303] = 6'd30;
    assign memory[2304] = 6'd29;
    assign memory[2305] = 6'd30;
    assign memory[2306] = 6'd31;
    assign memory[2307] = 6'd31;
    assign memory[2308] = 6'd30;
    assign memory[2309] = 6'd30;
    assign memory[2310] = 6'd30;
    assign memory[2311] = 6'd30;
    assign memory[2312] = 6'd30;
    assign memory[2313] = 6'd30;
    assign memory[2314] = 6'd31;
    assign memory[2315] = 6'd31;
    assign memory[2316] = 6'd30;
    assign memory[2317] = 6'd30;
    assign memory[2318] = 6'd30;
    assign memory[2319] = 6'd31;
    assign memory[2320] = 6'd30;
    assign memory[2321] = 6'd30;
    assign memory[2322] = 6'd30;
    assign memory[2323] = 6'd30;
    assign memory[2324] = 6'd30;
    assign memory[2325] = 6'd29;
    assign memory[2326] = 6'd29;
    assign memory[2327] = 6'd30;
    assign memory[2328] = 6'd30;
    assign memory[2329] = 6'd30;
    assign memory[2330] = 6'd32;
    assign memory[2331] = 6'd34;
    assign memory[2332] = 6'd34;
    assign memory[2333] = 6'd32;
    assign memory[2334] = 6'd30;
    assign memory[2335] = 6'd30;
    assign memory[2336] = 6'd30;
    assign memory[2337] = 6'd31;
    assign memory[2338] = 6'd30;
    assign memory[2339] = 6'd32;
    assign memory[2340] = 6'd34;
    assign memory[2341] = 6'd33;
    assign memory[2342] = 6'd33;
    assign memory[2343] = 6'd33;
    assign memory[2344] = 6'd33;
    assign memory[2345] = 6'd33;
    assign memory[2346] = 6'd31;
    assign memory[2347] = 6'd31;
    assign memory[2348] = 6'd30;
    assign memory[2349] = 6'd30;
    assign memory[2350] = 6'd30;
    assign memory[2351] = 6'd31;
    assign memory[2352] = 6'd34;
    assign memory[2353] = 6'd34;
    assign memory[2354] = 6'd33;
    assign memory[2355] = 6'd31;
    assign memory[2356] = 6'd30;
    assign memory[2357] = 6'd31;
    assign memory[2358] = 6'd34;
    assign memory[2359] = 6'd33;
    assign memory[2360] = 6'd33;
    assign memory[2361] = 6'd33;
    assign memory[2362] = 6'd34;
    assign memory[2363] = 6'd33;
    assign memory[2364] = 6'd31;
    assign memory[2365] = 6'd29;
    assign memory[2366] = 6'd31;
    assign memory[2367] = 6'd33;
    assign memory[2368] = 6'd34;
    assign memory[2369] = 6'd33;
    assign memory[2370] = 6'd34;
    assign memory[2371] = 6'd34;
    assign memory[2372] = 6'd33;
    assign memory[2373] = 6'd33;
    assign memory[2374] = 6'd33;
    assign memory[2375] = 6'd32;
    assign memory[2376] = 6'd30;
    assign memory[2377] = 6'd29;
    assign memory[2378] = 6'd31;
    assign memory[2379] = 6'd33;
    assign memory[2380] = 6'd34;
    assign memory[2381] = 6'd34;
    assign memory[2382] = 6'd33;
    assign memory[2383] = 6'd33;
    assign memory[2384] = 6'd33;
    assign memory[2385] = 6'd34;
    assign memory[2386] = 6'd34;
    assign memory[2387] = 6'd33;
    assign memory[2388] = 6'd30;
    assign memory[2389] = 6'd30;
    assign memory[2390] = 6'd31;
    assign memory[2391] = 6'd33;
    assign memory[2392] = 6'd33;
    assign memory[2393] = 6'd33;
    assign memory[2394] = 6'd34;
    assign memory[2395] = 6'd34;
    assign memory[2396] = 6'd34;
    assign memory[2397] = 6'd33;
    assign memory[2398] = 6'd33;
    assign memory[2399] = 6'd32;
    assign memory[2400] = 6'd30;
    assign memory[2401] = 6'd30;
    assign memory[2402] = 6'd31;
    assign memory[2403] = 6'd30;
    assign memory[2404] = 6'd30;
    assign memory[2405] = 6'd31;
    assign memory[2406] = 6'd30;
    assign memory[2407] = 6'd30;
    assign memory[2408] = 6'd29;
    assign memory[2409] = 6'd30;
    assign memory[2410] = 6'd30;
    assign memory[2411] = 6'd30;
    assign memory[2412] = 6'd31;
    assign memory[2413] = 6'd30;
    assign memory[2414] = 6'd32;
    assign memory[2415] = 6'd34;
    assign memory[2416] = 6'd34;
    assign memory[2417] = 6'd32;
    assign memory[2418] = 6'd29;
    assign memory[2419] = 6'd30;
    assign memory[2420] = 6'd31;
    assign memory[2421] = 6'd31;
    assign memory[2422] = 6'd31;
    assign memory[2423] = 6'd30;
    assign memory[2424] = 6'd30;
    assign memory[2425] = 6'd30;
    assign memory[2426] = 6'd30;
    assign memory[2427] = 6'd30;
    assign memory[2428] = 6'd30;
    assign memory[2429] = 6'd30;
    assign memory[2430] = 6'd30;
    assign memory[2431] = 6'd31;
    assign memory[2432] = 6'd31;
    assign memory[2433] = 6'd31;
    assign memory[2434] = 6'd30;
    assign memory[2435] = 6'd30;
    assign memory[2436] = 6'd31;
    assign memory[2437] = 6'd30;
    assign memory[2438] = 6'd30;
    assign memory[2439] = 6'd30;
    assign memory[2440] = 6'd30;
    assign memory[2441] = 6'd30;
    assign memory[2442] = 6'd30;
    assign memory[2443] = 6'd30;
    assign memory[2444] = 6'd31;
    assign memory[2445] = 6'd31;
    assign memory[2446] = 6'd31;
    assign memory[2447] = 6'd31;
    assign memory[2448] = 6'd33;
    assign memory[2449] = 6'd34;
    assign memory[2450] = 6'd33;
    assign memory[2451] = 6'd31;
    assign memory[2452] = 6'd30;
    assign memory[2453] = 6'd31;
    assign memory[2454] = 6'd30;
    assign memory[2455] = 6'd30;
    assign memory[2456] = 6'd31;
    assign memory[2457] = 6'd33;
    assign memory[2458] = 6'd34;
    assign memory[2459] = 6'd34;
    assign memory[2460] = 6'd34;
    assign memory[2461] = 6'd33;
    assign memory[2462] = 6'd34;
    assign memory[2463] = 6'd34;
    assign memory[2464] = 6'd34;
    assign memory[2465] = 6'd34;
    assign memory[2466] = 6'd34;
    assign memory[2467] = 6'd33;
    assign memory[2468] = 6'd33;
    assign memory[2469] = 6'd33;
    assign memory[2470] = 6'd33;
    assign memory[2471] = 6'd33;
    assign memory[2472] = 6'd33;
    assign memory[2473] = 6'd34;
    assign memory[2474] = 6'd33;
    assign memory[2475] = 6'd31;
    assign memory[2476] = 6'd29;
    assign memory[2477] = 6'd31;
    assign memory[2478] = 6'd33;
    assign memory[2479] = 6'd33;
    assign memory[2480] = 6'd33;
    assign memory[2481] = 6'd33;
    assign memory[2482] = 6'd34;
    assign memory[2483] = 6'd34;
    assign memory[2484] = 6'd34;
    assign memory[2485] = 6'd33;
    assign memory[2486] = 6'd33;
    assign memory[2487] = 6'd33;
    assign memory[2488] = 6'd33;
    assign memory[2489] = 6'd34;
    assign memory[2490] = 6'd33;
    assign memory[2491] = 6'd33;
    assign memory[2492] = 6'd33;
    assign memory[2493] = 6'd33;
    assign memory[2494] = 6'd33;
    assign memory[2495] = 6'd33;
    assign memory[2496] = 6'd33;
    assign memory[2497] = 6'd33;
    assign memory[2498] = 6'd33;
    assign memory[2499] = 6'd33;
    assign memory[2500] = 6'd34;
    assign memory[2501] = 6'd34;
    assign memory[2502] = 6'd34;
    assign memory[2503] = 6'd34;
    assign memory[2504] = 6'd34;
    assign memory[2505] = 6'd34;
    assign memory[2506] = 6'd33;
    assign memory[2507] = 6'd33;
    assign memory[2508] = 6'd33;
    assign memory[2509] = 6'd34;
    assign memory[2510] = 6'd34;
    assign memory[2511] = 6'd33;
    assign memory[2512] = 6'd33;
    assign memory[2513] = 6'd33;
    assign memory[2514] = 6'd33;
    assign memory[2515] = 6'd34;
    assign memory[2516] = 6'd33;
    assign memory[2517] = 6'd31;
    assign memory[2518] = 6'd30;
    assign memory[2519] = 6'd31;
    assign memory[2520] = 6'd33;
    assign memory[2521] = 6'd34;
    assign memory[2522] = 6'd33;
    assign memory[2523] = 6'd34;
    assign memory[2524] = 6'd34;
    assign memory[2525] = 6'd33;
    assign memory[2526] = 6'd30;
    assign memory[2527] = 6'd30;
    assign memory[2528] = 6'd31;
    assign memory[2529] = 6'd33;
    assign memory[2530] = 6'd34;
    assign memory[2531] = 6'd34;
    assign memory[2532] = 6'd34;
    assign memory[2533] = 6'd34;
    assign memory[2534] = 6'd34;
    assign memory[2535] = 6'd31;
    assign memory[2536] = 6'd30;
    assign memory[2537] = 6'd30;
    assign memory[2538] = 6'd30;
    assign memory[2539] = 6'd29;
    assign memory[2540] = 6'd30;
    assign memory[2541] = 6'd33;
    assign memory[2542] = 6'd34;
    assign memory[2543] = 6'd33;
    assign memory[2544] = 6'd31;
    assign memory[2545] = 6'd30;
    assign memory[2546] = 6'd31;
    assign memory[2547] = 6'd30;
    assign memory[2548] = 6'd30;
    assign memory[2549] = 6'd31;
    assign memory[2550] = 6'd33;
    assign memory[2551] = 6'd34;
    assign memory[2552] = 6'd33;
    assign memory[2553] = 6'd30;
    assign memory[2554] = 6'd29;
    assign memory[2555] = 6'd31;
    assign memory[2556] = 6'd30;
    assign memory[2557] = 6'd31;
    assign memory[2558] = 6'd30;
    assign memory[2559] = 6'd30;
    assign memory[2560] = 6'd30;
    assign memory[2561] = 6'd30;
    assign memory[2562] = 6'd30;
    assign memory[2563] = 6'd30;
    assign memory[2564] = 6'd31;
    assign memory[2565] = 6'd31;
    assign memory[2566] = 6'd30;
    assign memory[2567] = 6'd31;
    assign memory[2568] = 6'd33;
    assign memory[2569] = 6'd34;
    assign memory[2570] = 6'd33;
    assign memory[2571] = 6'd31;
    assign memory[2572] = 6'd30;
    assign memory[2573] = 6'd31;
    assign memory[2574] = 6'd30;
    assign memory[2575] = 6'd30;
    assign memory[2576] = 6'd31;
    assign memory[2577] = 6'd31;
    assign memory[2578] = 6'd30;
    assign memory[2579] = 6'd30;
    assign memory[2580] = 6'd30;
    assign memory[2581] = 6'd31;
    assign memory[2582] = 6'd30;
    assign memory[2583] = 6'd30;
    assign memory[2584] = 6'd30;
    assign memory[2585] = 6'd30;
    assign memory[2586] = 6'd31;
    assign memory[2587] = 6'd31;
    assign memory[2588] = 6'd31;
    assign memory[2589] = 6'd30;
    assign memory[2590] = 6'd30;
    assign memory[2591] = 6'd30;
    assign memory[2592] = 6'd30;
    assign memory[2593] = 6'd30;
    assign memory[2594] = 6'd31;
    assign memory[2595] = 6'd31;
    assign memory[2596] = 6'd30;
    assign memory[2597] = 6'd31;
    assign memory[2598] = 6'd33;
    assign memory[2599] = 6'd34;
    assign memory[2600] = 6'd33;
    assign memory[2601] = 6'd31;
    assign memory[2602] = 6'd30;
    assign memory[2603] = 6'd31;
    assign memory[2604] = 6'd31;
    assign memory[2605] = 6'd30;
    assign memory[2606] = 6'd31;
    assign memory[2607] = 6'd32;
    assign memory[2608] = 6'd34;
    assign memory[2609] = 6'd33;
    assign memory[2610] = 6'd31;
    assign memory[2611] = 6'd30;
    assign memory[2612] = 6'd31;
    assign memory[2613] = 6'd33;
    assign memory[2614] = 6'd34;
    assign memory[2615] = 6'd33;
    assign memory[2616] = 6'd31;
    assign memory[2617] = 6'd30;
    assign memory[2618] = 6'd31;
    assign memory[2619] = 6'd30;
    assign memory[2620] = 6'd30;
    assign memory[2621] = 6'd30;
    assign memory[2622] = 6'd30;
    assign memory[2623] = 6'd30;
    assign memory[2624] = 6'd31;
    assign memory[2625] = 6'd33;
    assign memory[2626] = 6'd34;
    assign memory[2627] = 6'd33;
    assign memory[2628] = 6'd31;
    assign memory[2629] = 6'd30;
    assign memory[2630] = 6'd31;
    assign memory[2631] = 6'd32;
    assign memory[2632] = 6'd33;
    assign memory[2633] = 6'd32;
    assign memory[2634] = 6'd33;
    assign memory[2635] = 6'd32;
    assign memory[2636] = 6'd33;
    assign memory[2637] = 6'd34;
    assign memory[2638] = 6'd33;
    assign memory[2639] = 6'd33;
    assign memory[2640] = 6'd33;
    assign memory[2641] = 6'd33;
    assign memory[2642] = 6'd34;
    assign memory[2643] = 6'd34;
    assign memory[2644] = 6'd34;
    assign memory[2645] = 6'd33;
    assign memory[2646] = 6'd33;
    assign memory[2647] = 6'd33;
    assign memory[2648] = 6'd33;
    assign memory[2649] = 6'd33;
    assign memory[2650] = 6'd33;
    assign memory[2651] = 6'd33;
    assign memory[2652] = 6'd33;
    assign memory[2653] = 6'd33;
    assign memory[2654] = 6'd33;
    assign memory[2655] = 6'd31;
    assign memory[2656] = 6'd29;
    assign memory[2657] = 6'd30;
    assign memory[2658] = 6'd30;
    assign memory[2659] = 6'd30;
    assign memory[2660] = 6'd30;
    assign memory[2661] = 6'd33;
    assign memory[2662] = 6'd34;
    assign memory[2663] = 6'd33;
    assign memory[2664] = 6'd33;
    assign memory[2665] = 6'd34;
    assign memory[2666] = 6'd34;
    assign memory[2667] = 6'd34;
    assign memory[2668] = 6'd34;
    assign memory[2669] = 6'd33;
    assign memory[2670] = 6'd33;
    assign memory[2671] = 6'd33;
    assign memory[2672] = 6'd34;
    assign memory[2673] = 6'd34;
    assign memory[2674] = 6'd33;
    assign memory[2675] = 6'd34;
    assign memory[2676] = 6'd34;
    assign memory[2677] = 6'd33;
    assign memory[2678] = 6'd33;
    assign memory[2679] = 6'd34;
    assign memory[2680] = 6'd33;
    assign memory[2681] = 6'd34;
    assign memory[2682] = 6'd33;
    assign memory[2683] = 6'd33;
    assign memory[2684] = 6'd33;
    assign memory[2685] = 6'd34;
    assign memory[2686] = 6'd33;
    assign memory[2687] = 6'd34;
    assign memory[2688] = 6'd33;
    assign memory[2689] = 6'd34;
    assign memory[2690] = 6'd33;
    assign memory[2691] = 6'd33;
    assign memory[2692] = 6'd34;
    assign memory[2693] = 6'd34;
    assign memory[2694] = 6'd33;
    assign memory[2695] = 6'd34;
    assign memory[2696] = 6'd34;
    assign memory[2697] = 6'd32;
    assign memory[2698] = 6'd30;
    assign memory[2699] = 6'd31;
    assign memory[2700] = 6'd33;
    assign memory[2701] = 6'd34;
    assign memory[2702] = 6'd33;
    assign memory[2703] = 6'd34;
    assign memory[2704] = 6'd33;
    assign memory[2705] = 6'd33;
    assign memory[2706] = 6'd33;
    assign memory[2707] = 6'd34;
    assign memory[2708] = 6'd34;
    assign memory[2709] = 6'd31;
    assign memory[2710] = 6'd31;
    assign memory[2711] = 6'd31;
    assign memory[2712] = 6'd30;
    assign memory[2713] = 6'd31;
    assign memory[2714] = 6'd31;
    assign memory[2715] = 6'd33;
    assign memory[2716] = 6'd34;
    assign memory[2717] = 6'd34;
    assign memory[2718] = 6'd32;
    assign memory[2719] = 6'd31;
    assign memory[2720] = 6'd31;
    assign memory[2721] = 6'd30;
    assign memory[2722] = 6'd30;
    assign memory[2723] = 6'd30;
    assign memory[2724] = 6'd30;
    assign memory[2725] = 6'd31;
    assign memory[2726] = 6'd31;
    assign memory[2727] = 6'd31;
    assign memory[2728] = 6'd31;
    assign memory[2729] = 6'd31;
    assign memory[2730] = 6'd31;
    assign memory[2731] = 6'd30;
    assign memory[2732] = 6'd30;
    assign memory[2733] = 6'd29;
    assign memory[2734] = 6'd30;
    assign memory[2735] = 6'd30;
    assign memory[2736] = 6'd30;
    assign memory[2737] = 6'd29;
    assign memory[2738] = 6'd30;
    assign memory[2739] = 6'd31;
    assign memory[2740] = 6'd30;
    assign memory[2741] = 6'd30;
    assign memory[2742] = 6'd30;
    assign memory[2743] = 6'd30;
    assign memory[2744] = 6'd30;
    assign memory[2745] = 6'd30;
    assign memory[2746] = 6'd29;
    assign memory[2747] = 6'd30;
    assign memory[2748] = 6'd30;
    assign memory[2749] = 6'd30;
    assign memory[2750] = 6'd30;
    assign memory[2751] = 6'd33;
    assign memory[2752] = 6'd34;
    assign memory[2753] = 6'd34;
    assign memory[2754] = 6'd31;
    assign memory[2755] = 6'd30;
    assign memory[2756] = 6'd30;
    assign memory[2757] = 6'd32;
    assign memory[2758] = 6'd34;
    assign memory[2759] = 6'd34;
    assign memory[2760] = 6'd31;
    assign memory[2761] = 6'd30;
    assign memory[2762] = 6'd30;
    assign memory[2763] = 6'd30;
    assign memory[2764] = 6'd30;
    assign memory[2765] = 6'd31;
    assign memory[2766] = 6'd30;
    assign memory[2767] = 6'd29;
    assign memory[2768] = 6'd30;
    assign memory[2769] = 6'd32;
    assign memory[2770] = 6'd34;
    assign memory[2771] = 6'd34;
    assign memory[2772] = 6'd31;
    assign memory[2773] = 6'd30;
    assign memory[2774] = 6'd30;
    assign memory[2775] = 6'd30;
    assign memory[2776] = 6'd30;
    assign memory[2777] = 6'd30;
    assign memory[2778] = 6'd33;
    assign memory[2779] = 6'd34;
    assign memory[2780] = 6'd33;
    assign memory[2781] = 6'd31;
    assign memory[2782] = 6'd30;
    assign memory[2783] = 6'd30;
    assign memory[2784] = 6'd29;
    assign memory[2785] = 6'd30;
    assign memory[2786] = 6'd30;
    assign memory[2787] = 6'd30;
    assign memory[2788] = 6'd30;
    assign memory[2789] = 6'd30;
    assign memory[2790] = 6'd29;
    assign memory[2791] = 6'd30;
    assign memory[2792] = 6'd30;
    assign memory[2793] = 6'd30;
    assign memory[2794] = 6'd30;
    assign memory[2795] = 6'd30;
    assign memory[2796] = 6'd32;
    assign memory[2797] = 6'd33;
    assign memory[2798] = 6'd33;
    assign memory[2799] = 6'd31;
    assign memory[2800] = 6'd30;
    assign memory[2801] = 6'd30;
    assign memory[2802] = 6'd33;
    assign memory[2803] = 6'd34;
    assign memory[2804] = 6'd33;
    assign memory[2805] = 6'd33;
    assign memory[2806] = 6'd33;
    assign memory[2807] = 6'd33;
    assign memory[2808] = 6'd33;
    assign memory[2809] = 6'd33;
    assign memory[2810] = 6'd33;
    assign memory[2811] = 6'd33;
    assign memory[2812] = 6'd33;
    assign memory[2813] = 6'd33;
    assign memory[2814] = 6'd33;
    assign memory[2815] = 6'd33;
    assign memory[2816] = 6'd34;
    assign memory[2817] = 6'd33;
    assign memory[2818] = 6'd33;
    assign memory[2819] = 6'd33;
    assign memory[2820] = 6'd33;
    assign memory[2821] = 6'd33;
    assign memory[2822] = 6'd34;
    assign memory[2823] = 6'd34;
    assign memory[2824] = 6'd33;
    assign memory[2825] = 6'd33;
    assign memory[2826] = 6'd33;
    assign memory[2827] = 6'd33;
    assign memory[2828] = 6'd34;
    assign memory[2829] = 6'd34;
    assign memory[2830] = 6'd33;
    assign memory[2831] = 6'd33;
    assign memory[2832] = 6'd33;
    assign memory[2833] = 6'd33;
    assign memory[2834] = 6'd33;
    assign memory[2835] = 6'd33;
    assign memory[2836] = 6'd34;
    assign memory[2837] = 6'd34;
    assign memory[2838] = 6'd32;
    assign memory[2839] = 6'd30;
    assign memory[2840] = 6'd30;
    assign memory[2841] = 6'd30;
    assign memory[2842] = 6'd30;
    assign memory[2843] = 6'd30;
    assign memory[2844] = 6'd32;
    assign memory[2845] = 6'd34;
    assign memory[2846] = 6'd34;
    assign memory[2847] = 6'd30;
    assign memory[2848] = 6'd30;
    assign memory[2849] = 6'd31;
    assign memory[2850] = 6'd31;
    assign memory[2851] = 6'd31;
    assign memory[2852] = 6'd30;
    assign memory[2853] = 6'd30;
    assign memory[2854] = 6'd30;
    assign memory[2855] = 6'd30;
    assign memory[2856] = 6'd31;
    assign memory[2857] = 6'd30;
    assign memory[2858] = 6'd31;
    assign memory[2859] = 6'd33;
    assign memory[2860] = 6'd35;
    assign memory[2861] = 6'd34;
    assign memory[2862] = 6'd32;
    assign memory[2863] = 6'd30;
    assign memory[2864] = 6'd30;
    assign memory[2865] = 6'd30;
    assign memory[2866] = 6'd30;
    assign memory[2867] = 6'd31;
    assign memory[2868] = 6'd31;
    assign memory[2869] = 6'd30;
    assign memory[2870] = 6'd30;
    assign memory[2871] = 6'd31;
    assign memory[2872] = 6'd31;
    assign memory[2873] = 6'd31;
    assign memory[2874] = 6'd31;
    assign memory[2875] = 6'd31;
    assign memory[2876] = 6'd30;
    assign memory[2877] = 6'd31;
    assign memory[2878] = 6'd31;
    assign memory[2879] = 6'd31;
    assign memory[2880] = 6'd30;
    assign memory[2881] = 6'd30;
    assign memory[2882] = 6'd30;
    assign memory[2883] = 6'd30;
    assign memory[2884] = 6'd30;
    assign memory[2885] = 6'd30;
    assign memory[2886] = 6'd31;
    assign memory[2887] = 6'd31;
    assign memory[2888] = 6'd31;
    assign memory[2889] = 6'd33;
    assign memory[2890] = 6'd34;
    assign memory[2891] = 6'd33;
    assign memory[2892] = 6'd32;
    assign memory[2893] = 6'd30;
    assign memory[2894] = 6'd29;
    assign memory[2895] = 6'd30;
    assign memory[2896] = 6'd29;
    assign memory[2897] = 6'd30;
    assign memory[2898] = 6'd29;
    assign memory[2899] = 6'd31;
    assign memory[2900] = 6'd31;
    assign memory[2901] = 6'd32;
    assign memory[2902] = 6'd34;
    assign memory[2903] = 6'd34;
    assign memory[2904] = 6'd32;
    assign memory[2905] = 6'd31;
    assign memory[2906] = 6'd30;
    assign memory[2907] = 6'd31;
    assign memory[2908] = 6'd30;
    assign memory[2909] = 6'd30;
    assign memory[2910] = 6'd31;
    assign memory[2911] = 6'd30;
    assign memory[2912] = 6'd30;
    assign memory[2913] = 6'd32;
    assign memory[2914] = 6'd34;
    assign memory[2915] = 6'd33;
    assign memory[2916] = 6'd32;
    assign memory[2917] = 6'd30;
    assign memory[2918] = 6'd30;
    assign memory[2919] = 6'd32;
    assign memory[2920] = 6'd34;
    assign memory[2921] = 6'd33;
    assign memory[2922] = 6'd33;
    assign memory[2923] = 6'd34;
    assign memory[2924] = 6'd33;
    assign memory[2925] = 6'd32;
    assign memory[2926] = 6'd30;
    assign memory[2927] = 6'd30;
    assign memory[2928] = 6'd32;
    assign memory[2929] = 6'd33;
    assign memory[2930] = 6'd34;
    assign memory[2931] = 6'd34;
    assign memory[2932] = 6'd33;
    assign memory[2933] = 6'd33;
    assign memory[2934] = 6'd33;
    assign memory[2935] = 6'd33;
    assign memory[2936] = 6'd33;
    assign memory[2937] = 6'd32;
    assign memory[2938] = 6'd29;
    assign memory[2939] = 6'd30;
    assign memory[2940] = 6'd32;
    assign memory[2941] = 6'd33;
    assign memory[2942] = 6'd34;
    assign memory[2943] = 6'd33;
    assign memory[2944] = 6'd34;
    assign memory[2945] = 6'd33;
    assign memory[2946] = 6'd33;
    assign memory[2947] = 6'd33;
    assign memory[2948] = 6'd33;
    assign memory[2949] = 6'd33;
    assign memory[2950] = 6'd34;
    assign memory[2951] = 6'd34;
    assign memory[2952] = 6'd33;
    assign memory[2953] = 6'd33;
    assign memory[2954] = 6'd33;
    assign memory[2955] = 6'd33;
    assign memory[2956] = 6'd34;
    assign memory[2957] = 6'd33;
    assign memory[2958] = 6'd34;
    assign memory[2959] = 6'd34;
    assign memory[2960] = 6'd34;
    assign memory[2961] = 6'd34;
    assign memory[2962] = 6'd34;
    assign memory[2963] = 6'd34;
    assign memory[2964] = 6'd34;
    assign memory[2965] = 6'd33;
    assign memory[2966] = 6'd33;
    assign memory[2967] = 6'd33;
    assign memory[2968] = 6'd33;
    assign memory[2969] = 6'd34;
    assign memory[2970] = 6'd34;
    assign memory[2971] = 6'd34;
    assign memory[2972] = 6'd34;
    assign memory[2973] = 6'd34;
    assign memory[2974] = 6'd34;
    assign memory[2975] = 6'd34;
    assign memory[2976] = 6'd34;
    assign memory[2977] = 6'd33;
    assign memory[2978] = 6'd33;
    assign memory[2979] = 6'd33;
    assign memory[2980] = 6'd33;
    assign memory[2981] = 6'd34;
    assign memory[2982] = 6'd31;
    assign memory[2983] = 6'd30;
    assign memory[2984] = 6'd30;
    assign memory[2985] = 6'd31;
    assign memory[2986] = 6'd30;
    assign memory[2987] = 6'd30;
    assign memory[2988] = 6'd30;
    assign memory[2989] = 6'd30;
    assign memory[2990] = 6'd30;
    assign memory[2991] = 6'd30;
    assign memory[2992] = 6'd31;
    assign memory[2993] = 6'd30;
    assign memory[2994] = 6'd30;
    assign memory[2995] = 6'd30;
    assign memory[2996] = 6'd30;
    assign memory[2997] = 6'd30;
    assign memory[2998] = 6'd30;
    assign memory[2999] = 6'd30;
    assign memory[3000] = 6'd31;
    assign memory[3001] = 6'd31;
    assign memory[3002] = 6'd31;
    assign memory[3003] = 6'd31;
    assign memory[3004] = 6'd30;
    assign memory[3005] = 6'd30;
    assign memory[3006] = 6'd29;
    assign memory[3007] = 6'd29;
    assign memory[3008] = 6'd30;
    assign memory[3009] = 6'd30;
    assign memory[3010] = 6'd30;
    assign memory[3011] = 6'd30;
    assign memory[3012] = 6'd31;
    assign memory[3013] = 6'd31;
    assign memory[3014] = 6'd30;
    assign memory[3015] = 6'd30;
    assign memory[3016] = 6'd31;
    assign memory[3017] = 6'd30;
    assign memory[3018] = 6'd30;
    assign memory[3019] = 6'd30;
    assign memory[3020] = 6'd30;
    assign memory[3021] = 6'd30;
    assign memory[3022] = 6'd30;
    assign memory[3023] = 6'd30;
    assign memory[3024] = 6'd30;
    assign memory[3025] = 6'd30;
    assign memory[3026] = 6'd30;
    assign memory[3027] = 6'd31;
    assign memory[3028] = 6'd31;
    assign memory[3029] = 6'd31;
    assign memory[3030] = 6'd30;
    assign memory[3031] = 6'd30;
    assign memory[3032] = 6'd31;
    assign memory[3033] = 6'd31;
    assign memory[3034] = 6'd31;
    assign memory[3035] = 6'd31;
    assign memory[3036] = 6'd30;
    assign memory[3037] = 6'd30;
    assign memory[3038] = 6'd30;
    assign memory[3039] = 6'd30;
    assign memory[3040] = 6'd30;
    assign memory[3041] = 6'd30;
    assign memory[3042] = 6'd32;
    assign memory[3043] = 6'd34;
    assign memory[3044] = 6'd34;
    assign memory[3045] = 6'd32;
    assign memory[3046] = 6'd31;
    assign memory[3047] = 6'd31;
    assign memory[3048] = 6'd30;
    assign memory[3049] = 6'd30;
    assign memory[3050] = 6'd31;
    assign memory[3051] = 6'd32;
    assign memory[3052] = 6'd34;
    assign memory[3053] = 6'd34;
    assign memory[3054] = 6'd34;
    assign memory[3055] = 6'd33;
    assign memory[3056] = 6'd33;
    assign memory[3057] = 6'd32;
    assign memory[3058] = 6'd30;
    assign memory[3059] = 6'd31;
    assign memory[3060] = 6'd30;
    assign memory[3061] = 6'd31;
    assign memory[3062] = 6'd30;
    assign memory[3063] = 6'd30;
    assign memory[3064] = 6'd30;
    assign memory[3065] = 6'd30;
    assign memory[3066] = 6'd32;
    assign memory[3067] = 6'd33;
    assign memory[3068] = 6'd34;
    assign memory[3069] = 6'd31;
    assign memory[3070] = 6'd30;
    assign memory[3071] = 6'd30;
    assign memory[3072] = 6'd32;
    assign memory[3073] = 6'd33;
    assign memory[3074] = 6'd34;
    assign memory[3075] = 6'd32;
    assign memory[3076] = 6'd30;
    assign memory[3077] = 6'd30;
    assign memory[3078] = 6'd31;
    assign memory[3079] = 6'd30;
    assign memory[3080] = 6'd30;
    assign memory[3081] = 6'd30;
    assign memory[3082] = 6'd30;
    assign memory[3083] = 6'd30;
    assign memory[3084] = 6'd31;
    assign memory[3085] = 6'd30;
    assign memory[3086] = 6'd31;
    assign memory[3087] = 6'd30;
    assign memory[3088] = 6'd30;
    assign memory[3089] = 6'd30;
    assign memory[3090] = 6'd31;
    assign memory[3091] = 6'd30;
    assign memory[3092] = 6'd30;
    assign memory[3093] = 6'd30;
    assign memory[3094] = 6'd29;
    assign memory[3095] = 6'd30;
    assign memory[3096] = 6'd30;
    assign memory[3097] = 6'd30;
    assign memory[3098] = 6'd31;
    assign memory[3099] = 6'd31;
    assign memory[3100] = 6'd30;
    assign memory[3101] = 6'd30;
    assign memory[3102] = 6'd30;
    assign memory[3103] = 6'd30;
    assign memory[3104] = 6'd30;
    assign memory[3105] = 6'd30;
    assign memory[3106] = 6'd30;
    assign memory[3107] = 6'd30;
    assign memory[3108] = 6'd30;
    assign memory[3109] = 6'd30;
    assign memory[3110] = 6'd30;
    assign memory[3111] = 6'd30;
    assign memory[3112] = 6'd30;
    assign memory[3113] = 6'd29;
    assign memory[3114] = 6'd30;
    assign memory[3115] = 6'd30;
    assign memory[3116] = 6'd31;
    assign memory[3117] = 6'd30;
    assign memory[3118] = 6'd30;
    assign memory[3119] = 6'd30;
    assign memory[3120] = 6'd30;
    assign memory[3121] = 6'd30;
    assign memory[3122] = 6'd29;
    assign memory[3123] = 6'd30;
    assign memory[3124] = 6'd31;
    assign memory[3125] = 6'd30;
    assign memory[3126] = 6'd30;
    assign memory[3127] = 6'd31;
    assign memory[3128] = 6'd30;
    assign memory[3129] = 6'd30;
    assign memory[3130] = 6'd30;
    assign memory[3131] = 6'd30;
    assign memory[3132] = 6'd30;
    assign memory[3133] = 6'd30;
    assign memory[3134] = 6'd30;
    assign memory[3135] = 6'd31;
    assign memory[3136] = 6'd31;
    assign memory[3137] = 6'd30;
    assign memory[3138] = 6'd30;
    assign memory[3139] = 6'd30;
    assign memory[3140] = 6'd30;
    assign memory[3141] = 6'd30;
    assign memory[3142] = 6'd30;
    assign memory[3143] = 6'd30;
    assign memory[3144] = 6'd30;
    assign memory[3145] = 6'd30;
    assign memory[3146] = 6'd30;
    assign memory[3147] = 6'd30;
    assign memory[3148] = 6'd30;
    assign memory[3149] = 6'd30;
    assign memory[3150] = 6'd31;
    assign memory[3151] = 6'd30;
    assign memory[3152] = 6'd30;
    assign memory[3153] = 6'd31;
    assign memory[3154] = 6'd30;
    assign memory[3155] = 6'd29;
    assign memory[3156] = 6'd30;
    assign memory[3157] = 6'd30;
    assign memory[3158] = 6'd31;
    assign memory[3159] = 6'd31;
    assign memory[3160] = 6'd30;
    assign memory[3161] = 6'd30;
    assign memory[3162] = 6'd30;
    assign memory[3163] = 6'd30;
    assign memory[3164] = 6'd30;
    assign memory[3165] = 6'd30;
    assign memory[3166] = 6'd30;
    assign memory[3167] = 6'd31;
    assign memory[3168] = 6'd31;
    assign memory[3169] = 6'd30;
    assign memory[3170] = 6'd30;
    assign memory[3171] = 6'd30;
    assign memory[3172] = 6'd30;
    assign memory[3173] = 6'd31;
    assign memory[3174] = 6'd31;
    assign memory[3175] = 6'd30;
    assign memory[3176] = 6'd31;
    assign memory[3177] = 6'd31;
    assign memory[3178] = 6'd30;
    assign memory[3179] = 6'd30;
    assign memory[3180] = 6'd30;
    assign memory[3181] = 6'd30;
    assign memory[3182] = 6'd31;
    assign memory[3183] = 6'd31;
    assign memory[3184] = 6'd31;
    assign memory[3185] = 6'd31;
    assign memory[3186] = 6'd30;
    assign memory[3187] = 6'd31;
    assign memory[3188] = 6'd30;
    assign memory[3189] = 6'd31;
    assign memory[3190] = 6'd30;
    assign memory[3191] = 6'd31;
    assign memory[3192] = 6'd31;
    assign memory[3193] = 6'd31;
    assign memory[3194] = 6'd31;
    assign memory[3195] = 6'd31;
    assign memory[3196] = 6'd30;
    assign memory[3197] = 6'd30;
    assign memory[3198] = 6'd30;
    assign memory[3199] = 6'd31;
    assign memory[3200] = 6'd30;
    assign memory[3201] = 6'd30;
    assign memory[3202] = 6'd31;
    assign memory[3203] = 6'd30;
    assign memory[3204] = 6'd31;
    assign memory[3205] = 6'd30;
    assign memory[3206] = 6'd30;
    assign memory[3207] = 6'd29;
    assign memory[3208] = 6'd30;
    assign memory[3209] = 6'd30;
    assign memory[3210] = 6'd30;
    assign memory[3211] = 6'd30;
    assign memory[3212] = 6'd30;
    assign memory[3213] = 6'd30;
    assign memory[3214] = 6'd30;
    assign memory[3215] = 6'd30;
    assign memory[3216] = 6'd31;
    assign memory[3217] = 6'd30;
    assign memory[3218] = 6'd30;
    assign memory[3219] = 6'd30;
    assign memory[3220] = 6'd30;
    assign memory[3221] = 6'd30;
    assign memory[3222] = 6'd30;
    assign memory[3223] = 6'd30;
    assign memory[3224] = 6'd30;
    assign memory[3225] = 6'd31;
    assign memory[3226] = 6'd30;
    assign memory[3227] = 6'd30;
    assign memory[3228] = 6'd30;
    assign memory[3229] = 6'd30;
    assign memory[3230] = 6'd30;
    assign memory[3231] = 6'd30;
    assign memory[3232] = 6'd30;
    assign memory[3233] = 6'd30;
    assign memory[3234] = 6'd30;
    assign memory[3235] = 6'd30;
    assign memory[3236] = 6'd32;
    assign memory[3237] = 6'd32;
    assign memory[3238] = 6'd32;
    assign memory[3239] = 6'd32;
    assign memory[3240] = 6'd32;
    assign memory[3241] = 6'd32;
    assign memory[3242] = 6'd31;
    assign memory[3243] = 6'd32;
    assign memory[3244] = 6'd31;
    assign memory[3245] = 6'd32;
    assign memory[3246] = 6'd31;
    assign memory[3247] = 6'd32;
    assign memory[3248] = 6'd32;
    assign memory[3249] = 6'd32;
    assign memory[3250] = 6'd32;
    assign memory[3251] = 6'd32;
    assign memory[3252] = 6'd32;
    assign memory[3253] = 6'd32;
    assign memory[3254] = 6'd32;
    assign memory[3255] = 6'd32;
    assign memory[3256] = 6'd32;
    assign memory[3257] = 6'd32;
    assign memory[3258] = 6'd32;
    assign memory[3259] = 6'd31;
    assign memory[3260] = 6'd32;
    assign memory[3261] = 6'd32;
    assign memory[3262] = 6'd32;
    assign memory[3263] = 6'd32;
    assign memory[3264] = 6'd31;
    assign memory[3265] = 6'd31;
    assign memory[3266] = 6'd32;
    assign memory[3267] = 6'd31;
    assign memory[3268] = 6'd32;
    assign memory[3269] = 6'd32;
    assign memory[3270] = 6'd32;
    assign memory[3271] = 6'd31;
    assign memory[3272] = 6'd32;
    assign memory[3273] = 6'd31;
    assign memory[3274] = 6'd31;
    assign memory[3275] = 6'd32;
    assign memory[3276] = 6'd31;
    assign memory[3277] = 6'd32;
    assign memory[3278] = 6'd32;
    assign memory[3279] = 6'd32;
    assign memory[3280] = 6'd32;
    assign memory[3281] = 6'd32;
    assign memory[3282] = 6'd32;
    assign memory[3283] = 6'd31;
    assign memory[3284] = 6'd32;
    assign memory[3285] = 6'd32;
    assign memory[3286] = 6'd32;
    assign memory[3287] = 6'd32;
    assign memory[3288] = 6'd31;
    assign memory[3289] = 6'd31;
    assign memory[3290] = 6'd31;
    assign memory[3291] = 6'd31;
    assign memory[3292] = 6'd32;
    assign memory[3293] = 6'd32;
    assign memory[3294] = 6'd32;
    assign memory[3295] = 6'd32;
    assign memory[3296] = 6'd31;
    assign memory[3297] = 6'd31;
    assign memory[3298] = 6'd32;
    assign memory[3299] = 6'd32;
    assign memory[3300] = 6'd32;
    assign memory[3301] = 6'd32;
    assign memory[3302] = 6'd32;
    assign memory[3303] = 6'd32;
    assign memory[3304] = 6'd32;
    assign memory[3305] = 6'd31;
    assign memory[3306] = 6'd32;
    assign memory[3307] = 6'd32;
    assign memory[3308] = 6'd31;
    assign memory[3309] = 6'd31;
    assign memory[3310] = 6'd31;
    assign memory[3311] = 6'd31;
    assign memory[3312] = 6'd32;
    assign memory[3313] = 6'd32;
    assign memory[3314] = 6'd32;
    assign memory[3315] = 6'd32;
    assign memory[3316] = 6'd32;
    assign memory[3317] = 6'd32;
    assign memory[3318] = 6'd32;
    assign memory[3319] = 6'd32;
    assign memory[3320] = 6'd32;
    assign memory[3321] = 6'd31;
    assign memory[3322] = 6'd32;
    assign memory[3323] = 6'd31;
    assign memory[3324] = 6'd32;
    assign memory[3325] = 6'd32;
    assign memory[3326] = 6'd32;
    assign memory[3327] = 6'd32;
    assign memory[3328] = 6'd32;
    assign memory[3329] = 6'd32;
    assign memory[3330] = 6'd32;
    assign memory[3331] = 6'd32;
    assign memory[3332] = 6'd32;
    assign memory[3333] = 6'd31;
    assign memory[3334] = 6'd32;
    assign memory[3335] = 6'd32;
    assign memory[3336] = 6'd32;
    assign memory[3337] = 6'd32;
    assign memory[3338] = 6'd32;
    assign memory[3339] = 6'd32;
    assign memory[3340] = 6'd32;
    assign memory[3341] = 6'd32;
    assign memory[3342] = 6'd32;
    assign memory[3343] = 6'd32;
    assign memory[3344] = 6'd32;
    assign memory[3345] = 6'd32;
    assign memory[3346] = 6'd32;
    assign memory[3347] = 6'd32;
    assign memory[3348] = 6'd32;
    assign memory[3349] = 6'd31;
    assign memory[3350] = 6'd32;
    assign memory[3351] = 6'd32;
    assign memory[3352] = 6'd32;
    assign memory[3353] = 6'd32;
    assign memory[3354] = 6'd32;
    assign memory[3355] = 6'd32;
    assign memory[3356] = 6'd32;
    assign memory[3357] = 6'd32;
    assign memory[3358] = 6'd31;
    assign memory[3359] = 6'd32;
    assign memory[3360] = 6'd31;
    assign memory[3361] = 6'd32;
    assign memory[3362] = 6'd32;
    assign memory[3363] = 6'd32;
    assign memory[3364] = 6'd32;
    assign memory[3365] = 6'd32;
    assign memory[3366] = 6'd32;
    assign memory[3367] = 6'd32;
    assign memory[3368] = 6'd31;
    assign memory[3369] = 6'd31;
    assign memory[3370] = 6'd32;
    assign memory[3371] = 6'd32;
    assign memory[3372] = 6'd32;
    assign memory[3373] = 6'd32;
    assign memory[3374] = 6'd31;
    assign memory[3375] = 6'd31;
    assign memory[3376] = 6'd31;
    assign memory[3377] = 6'd31;
    assign memory[3378] = 6'd32;
    assign memory[3379] = 6'd32;
    assign memory[3380] = 6'd32;
    assign memory[3381] = 6'd31;
    assign memory[3382] = 6'd32;
    assign memory[3383] = 6'd32;
    assign memory[3384] = 6'd32;
    assign memory[3385] = 6'd32;
    assign memory[3386] = 6'd32;
    assign memory[3387] = 6'd32;
    assign memory[3388] = 6'd32;
    assign memory[3389] = 6'd32;
    assign memory[3390] = 6'd32;
    assign memory[3391] = 6'd32;
    assign memory[3392] = 6'd32;
    assign memory[3393] = 6'd32;
    assign memory[3394] = 6'd31;
    assign memory[3395] = 6'd31;
    assign memory[3396] = 6'd32;
    assign memory[3397] = 6'd32;
    assign memory[3398] = 6'd31;
    assign memory[3399] = 6'd31;
    assign memory[3400] = 6'd32;
    assign memory[3401] = 6'd32;
    assign memory[3402] = 6'd31;
    assign memory[3403] = 6'd32;
    assign memory[3404] = 6'd33;
    assign memory[3405] = 6'd33;
    assign memory[3406] = 6'd32;
    assign memory[3407] = 6'd31;
    assign memory[3408] = 6'd31;
    assign memory[3409] = 6'd32;
    assign memory[3410] = 6'd32;
    assign memory[3411] = 6'd32;
    assign memory[3412] = 6'd32;
    assign memory[3413] = 6'd31;
    assign memory[3414] = 6'd31;
    assign memory[3415] = 6'd32;
    assign memory[3416] = 6'd32;
    assign memory[3417] = 6'd31;
    assign memory[3418] = 6'd31;
    assign memory[3419] = 6'd32;
    assign memory[3420] = 6'd32;
    assign memory[3421] = 6'd32;
    assign memory[3422] = 6'd32;
    assign memory[3423] = 6'd32;
    assign memory[3424] = 6'd32;
    assign memory[3425] = 6'd32;
    assign memory[3426] = 6'd32;
    assign memory[3427] = 6'd32;
    assign memory[3428] = 6'd32;
    assign memory[3429] = 6'd32;
    assign memory[3430] = 6'd32;
    assign memory[3431] = 6'd32;
    assign memory[3432] = 6'd32;
    assign memory[3433] = 6'd32;
    assign memory[3434] = 6'd32;
    assign memory[3435] = 6'd32;
    assign memory[3436] = 6'd31;
    assign memory[3437] = 6'd32;
    assign memory[3438] = 6'd32;
    assign memory[3439] = 6'd32;
    assign memory[3440] = 6'd32;
    assign memory[3441] = 6'd31;
    assign memory[3442] = 6'd32;
    assign memory[3443] = 6'd32;
    assign memory[3444] = 6'd32;
    assign memory[3445] = 6'd31;
    assign memory[3446] = 6'd31;
    assign memory[3447] = 6'd31;
    assign memory[3448] = 6'd31;
    assign memory[3449] = 6'd32;
    assign memory[3450] = 6'd32;
    assign memory[3451] = 6'd31;
    assign memory[3452] = 6'd31;
    assign memory[3453] = 6'd32;
    assign memory[3454] = 6'd31;
    assign memory[3455] = 6'd31;
    assign memory[3456] = 6'd32;
    assign memory[3457] = 6'd31;
    assign memory[3458] = 6'd31;
    assign memory[3459] = 6'd32;
    assign memory[3460] = 6'd32;
    assign memory[3461] = 6'd31;
    assign memory[3462] = 6'd32;
    assign memory[3463] = 6'd31;
    assign memory[3464] = 6'd31;
    assign memory[3465] = 6'd32;
    assign memory[3466] = 6'd32;
    assign memory[3467] = 6'd32;
    assign memory[3468] = 6'd33;
    assign memory[3469] = 6'd32;
    assign memory[3470] = 6'd32;
    assign memory[3471] = 6'd31;
    assign memory[3472] = 6'd32;
    assign memory[3473] = 6'd32;
    assign memory[3474] = 6'd32;
    assign memory[3475] = 6'd32;
    assign memory[3476] = 6'd32;
    assign memory[3477] = 6'd33;
    assign memory[3478] = 6'd32;
    assign memory[3479] = 6'd32;
    assign memory[3480] = 6'd31;
    assign memory[3481] = 6'd32;
    assign memory[3482] = 6'd33;
    assign memory[3483] = 6'd32;
    assign memory[3484] = 6'd32;
    assign memory[3485] = 6'd32;
    assign memory[3486] = 6'd32;
    assign memory[3487] = 6'd31;
    assign memory[3488] = 6'd32;
    assign memory[3489] = 6'd32;
    assign memory[3490] = 6'd32;
    assign memory[3491] = 6'd32;
    assign memory[3492] = 6'd31;
    assign memory[3493] = 6'd32;
    assign memory[3494] = 6'd32;
    assign memory[3495] = 6'd32;
    assign memory[3496] = 6'd32;
    assign memory[3497] = 6'd32;
    assign memory[3498] = 6'd31;
    assign memory[3499] = 6'd32;
    assign memory[3500] = 6'd32;
    assign memory[3501] = 6'd32;
    assign memory[3502] = 6'd32;
    assign memory[3503] = 6'd32;
    assign memory[3504] = 6'd32;
    assign memory[3505] = 6'd32;
    assign memory[3506] = 6'd32;
    assign memory[3507] = 6'd32;
    assign memory[3508] = 6'd32;
    assign memory[3509] = 6'd31;
    assign memory[3510] = 6'd32;
    assign memory[3511] = 6'd31;
    assign memory[3512] = 6'd31;
    assign memory[3513] = 6'd31;
    assign memory[3514] = 6'd31;
    assign memory[3515] = 6'd32;
    assign memory[3516] = 6'd32;
    assign memory[3517] = 6'd32;
    assign memory[3518] = 6'd31;
    assign memory[3519] = 6'd31;
    assign memory[3520] = 6'd31;
    assign memory[3521] = 6'd31;
    assign memory[3522] = 6'd31;
    assign memory[3523] = 6'd32;
    assign memory[3524] = 6'd31;
    assign memory[3525] = 6'd32;
    assign memory[3526] = 6'd31;
    assign memory[3527] = 6'd31;
    assign memory[3528] = 6'd31;
    assign memory[3529] = 6'd32;
    assign memory[3530] = 6'd31;
    assign memory[3531] = 6'd31;
    assign memory[3532] = 6'd32;
    assign memory[3533] = 6'd32;
    assign memory[3534] = 6'd32;
    assign memory[3535] = 6'd32;
    assign memory[3536] = 6'd31;
    assign memory[3537] = 6'd31;
    assign memory[3538] = 6'd31;
    assign memory[3539] = 6'd32;
    assign memory[3540] = 6'd32;
    assign memory[3541] = 6'd32;
    assign memory[3542] = 6'd32;
    assign memory[3543] = 6'd32;
    assign memory[3544] = 6'd32;
    assign memory[3545] = 6'd32;
    assign memory[3546] = 6'd32;
    assign memory[3547] = 6'd31;
    assign memory[3548] = 6'd32;
    assign memory[3549] = 6'd32;
    assign memory[3550] = 6'd32;
    assign memory[3551] = 6'd31;
    assign memory[3552] = 6'd31;
    assign memory[3553] = 6'd31;
    assign memory[3554] = 6'd31;
    assign memory[3555] = 6'd31;
    assign memory[3556] = 6'd32;
    assign memory[3557] = 6'd32;
    assign memory[3558] = 6'd32;
    assign memory[3559] = 6'd32;
    assign memory[3560] = 6'd32;
    assign memory[3561] = 6'd31;
    assign memory[3562] = 6'd32;
    assign memory[3563] = 6'd32;
    assign memory[3564] = 6'd32;
    assign memory[3565] = 6'd32;
    assign memory[3566] = 6'd32;
    assign memory[3567] = 6'd32;
    assign memory[3568] = 6'd32;
    assign memory[3569] = 6'd32;
    assign memory[3570] = 6'd32;
    assign memory[3571] = 6'd31;
    assign memory[3572] = 6'd32;
    assign memory[3573] = 6'd32;
    assign memory[3574] = 6'd31;
    assign memory[3575] = 6'd32;
    assign memory[3576] = 6'd31;
    assign memory[3577] = 6'd32;
    assign memory[3578] = 6'd31;
    assign memory[3579] = 6'd32;
    assign memory[3580] = 6'd32;
    assign memory[3581] = 6'd33;
    assign memory[3582] = 6'd32;
    assign memory[3583] = 6'd32;
    assign memory[3584] = 6'd31;
    assign memory[3585] = 6'd32;
    assign memory[3586] = 6'd32;
    assign memory[3587] = 6'd32;
    assign memory[3588] = 6'd31;
    assign memory[3589] = 6'd32;
    assign memory[3590] = 6'd32;
    assign memory[3591] = 6'd32;
    assign memory[3592] = 6'd32;
    assign memory[3593] = 6'd32;
    assign memory[3594] = 6'd31;
    assign memory[3595] = 6'd32;
    assign memory[3596] = 6'd32;
    assign memory[3597] = 6'd32;
    assign memory[3598] = 6'd32;
    assign memory[3599] = 6'd32;
    assign memory[3600] = 6'd32;
    assign memory[3601] = 6'd32;
    assign memory[3602] = 6'd32;
    assign memory[3603] = 6'd32;
    assign memory[3604] = 6'd32;
    assign memory[3605] = 6'd32;
    assign memory[3606] = 6'd31;
    assign memory[3607] = 6'd32;
    assign memory[3608] = 6'd32;
    assign memory[3609] = 6'd32;
    assign memory[3610] = 6'd32;
    assign memory[3611] = 6'd32;
    assign memory[3612] = 6'd32;
    assign memory[3613] = 6'd32;
    assign memory[3614] = 6'd32;
    assign memory[3615] = 6'd32;
    assign memory[3616] = 6'd32;
    assign memory[3617] = 6'd32;
    assign memory[3618] = 6'd32;
    assign memory[3619] = 6'd31;
    assign memory[3620] = 6'd32;
    assign memory[3621] = 6'd31;
    assign memory[3622] = 6'd32;
    assign memory[3623] = 6'd31;
    assign memory[3624] = 6'd32;
    assign memory[3625] = 6'd32;
    assign memory[3626] = 6'd32;
    assign memory[3627] = 6'd31;
    assign memory[3628] = 6'd31;
    assign memory[3629] = 6'd32;
    assign memory[3630] = 6'd32;
    assign memory[3631] = 6'd32;
    assign memory[3632] = 6'd32;
    assign memory[3633] = 6'd32;
    assign memory[3634] = 6'd32;
    assign memory[3635] = 6'd31;
    assign memory[3636] = 6'd32;
    assign memory[3637] = 6'd32;
    assign memory[3638] = 6'd32;
    assign memory[3639] = 6'd32;
    assign memory[3640] = 6'd32;
    assign memory[3641] = 6'd32;
    assign memory[3642] = 6'd32;
    assign memory[3643] = 6'd32;
    assign memory[3644] = 6'd32;
    assign memory[3645] = 6'd31;
    assign memory[3646] = 6'd31;
    assign memory[3647] = 6'd31;
    assign memory[3648] = 6'd32;
    assign memory[3649] = 6'd32;
    assign memory[3650] = 6'd32;
    assign memory[3651] = 6'd32;
    assign memory[3652] = 6'd32;
    assign memory[3653] = 6'd31;
    assign memory[3654] = 6'd31;
    assign memory[3655] = 6'd32;
    assign memory[3656] = 6'd32;
    assign memory[3657] = 6'd32;
    assign memory[3658] = 6'd32;
    assign memory[3659] = 6'd32;
    assign memory[3660] = 6'd32;
    assign memory[3661] = 6'd31;
    assign memory[3662] = 6'd32;
    assign memory[3663] = 6'd32;
    assign memory[3664] = 6'd31;
    assign memory[3665] = 6'd32;
    assign memory[3666] = 6'd32;
    assign memory[3667] = 6'd32;
    assign memory[3668] = 6'd32;
    assign memory[3669] = 6'd32;
    assign memory[3670] = 6'd32;
    assign memory[3671] = 6'd32;
    assign memory[3672] = 6'd32;
    assign memory[3673] = 6'd32;
    assign memory[3674] = 6'd32;
    assign memory[3675] = 6'd32;
    assign memory[3676] = 6'd32;
    assign memory[3677] = 6'd32;
    assign memory[3678] = 6'd32;
    assign memory[3679] = 6'd32;
    assign memory[3680] = 6'd32;
    assign memory[3681] = 6'd32;
    assign memory[3682] = 6'd32;
    assign memory[3683] = 6'd32;
    assign memory[3684] = 6'd32;
    assign memory[3685] = 6'd32;
    assign memory[3686] = 6'd32;
    assign memory[3687] = 6'd32;
    assign memory[3688] = 6'd31;
    assign memory[3689] = 6'd32;
    assign memory[3690] = 6'd32;
    assign memory[3691] = 6'd32;
    assign memory[3692] = 6'd32;
    assign memory[3693] = 6'd32;
    assign memory[3694] = 6'd32;
    assign memory[3695] = 6'd32;
    assign memory[3696] = 6'd32;
    assign memory[3697] = 6'd32;
    assign memory[3698] = 6'd32;
    assign memory[3699] = 6'd31;
    assign memory[3700] = 6'd32;
    assign memory[3701] = 6'd32;
    assign memory[3702] = 6'd32;
    assign memory[3703] = 6'd32;
    assign memory[3704] = 6'd32;
    assign memory[3705] = 6'd32;
    assign memory[3706] = 6'd32;
    assign memory[3707] = 6'd32;
    assign memory[3708] = 6'd32;
    assign memory[3709] = 6'd31;
    assign memory[3710] = 6'd31;
    assign memory[3711] = 6'd31;
    assign memory[3712] = 6'd31;
    assign memory[3713] = 6'd31;
    assign memory[3714] = 6'd32;
    assign memory[3715] = 6'd32;
    assign memory[3716] = 6'd32;
    assign memory[3717] = 6'd32;
    assign memory[3718] = 6'd32;
    assign memory[3719] = 6'd32;
    assign memory[3720] = 6'd32;
    assign memory[3721] = 6'd32;
    assign memory[3722] = 6'd31;
    assign memory[3723] = 6'd32;
    assign memory[3724] = 6'd32;
    assign memory[3725] = 6'd32;
    assign memory[3726] = 6'd31;
    assign memory[3727] = 6'd31;
    assign memory[3728] = 6'd31;
    assign memory[3729] = 6'd31;
    assign memory[3730] = 6'd31;
    assign memory[3731] = 6'd32;
    assign memory[3732] = 6'd32;
    assign memory[3733] = 6'd31;
    assign memory[3734] = 6'd32;
    assign memory[3735] = 6'd31;
    assign memory[3736] = 6'd32;
    assign memory[3737] = 6'd32;
    assign memory[3738] = 6'd32;
    assign memory[3739] = 6'd32;
    assign memory[3740] = 6'd31;
    assign memory[3741] = 6'd31;
    assign memory[3742] = 6'd32;
    assign memory[3743] = 6'd32;
    assign memory[3744] = 6'd32;
    assign memory[3745] = 6'd32;
    assign memory[3746] = 6'd32;
    assign memory[3747] = 6'd32;
    assign memory[3748] = 6'd32;
    assign memory[3749] = 6'd32;
    assign memory[3750] = 6'd32;
    assign memory[3751] = 6'd32;
    assign memory[3752] = 6'd32;
    assign memory[3753] = 6'd31;
    assign memory[3754] = 6'd31;
    assign memory[3755] = 6'd32;
    assign memory[3756] = 6'd32;
    assign memory[3757] = 6'd32;
    assign memory[3758] = 6'd32;
    assign memory[3759] = 6'd32;
    assign memory[3760] = 6'd32;
    assign memory[3761] = 6'd32;
    assign memory[3762] = 6'd32;
    assign memory[3763] = 6'd32;
    assign memory[3764] = 6'd32;
    assign memory[3765] = 6'd32;
    assign memory[3766] = 6'd32;
    assign memory[3767] = 6'd33;
    assign memory[3768] = 6'd32;
    assign memory[3769] = 6'd32;
    assign memory[3770] = 6'd32;
    assign memory[3771] = 6'd32;
    assign memory[3772] = 6'd32;
    assign memory[3773] = 6'd32;
    assign memory[3774] = 6'd32;
    assign memory[3775] = 6'd32;
    assign memory[3776] = 6'd32;
    assign memory[3777] = 6'd32;
    assign memory[3778] = 6'd32;
    assign memory[3779] = 6'd32;
    assign memory[3780] = 6'd32;
    assign memory[3781] = 6'd32;
    assign memory[3782] = 6'd32;
    assign memory[3783] = 6'd31;
    assign memory[3784] = 6'd32;
    assign memory[3785] = 6'd32;
    assign memory[3786] = 6'd32;
    assign memory[3787] = 6'd32;
    assign memory[3788] = 6'd32;
    assign memory[3789] = 6'd32;
    assign memory[3790] = 6'd32;
    assign memory[3791] = 6'd32;
    assign memory[3792] = 6'd32;
    assign memory[3793] = 6'd32;
    assign memory[3794] = 6'd31;
    assign memory[3795] = 6'd32;
    assign memory[3796] = 6'd31;
    assign memory[3797] = 6'd32;
    assign memory[3798] = 6'd32;
    assign memory[3799] = 6'd31;
    assign memory[3800] = 6'd32;
    assign memory[3801] = 6'd32;
    assign memory[3802] = 6'd32;
    assign memory[3803] = 6'd31;
    assign memory[3804] = 6'd31;
    assign memory[3805] = 6'd31;
    assign memory[3806] = 6'd32;
    assign memory[3807] = 6'd31;
    assign memory[3808] = 6'd32;
    assign memory[3809] = 6'd32;
    assign memory[3810] = 6'd32;
    assign memory[3811] = 6'd32;
    assign memory[3812] = 6'd31;
    assign memory[3813] = 6'd32;
    assign memory[3814] = 6'd32;
    assign memory[3815] = 6'd32;
    assign memory[3816] = 6'd32;
    assign memory[3817] = 6'd31;
    assign memory[3818] = 6'd32;
    assign memory[3819] = 6'd32;
    assign memory[3820] = 6'd32;
    assign memory[3821] = 6'd32;
    assign memory[3822] = 6'd32;
    assign memory[3823] = 6'd32;
    assign memory[3824] = 6'd32;
    assign memory[3825] = 6'd32;
    assign memory[3826] = 6'd32;
    assign memory[3827] = 6'd31;
    assign memory[3828] = 6'd31;
    assign memory[3829] = 6'd32;
    assign memory[3830] = 6'd31;
    assign memory[3831] = 6'd32;
    assign memory[3832] = 6'd31;
    assign memory[3833] = 6'd32;
    assign memory[3834] = 6'd32;
    assign memory[3835] = 6'd31;
    assign memory[3836] = 6'd32;
    assign memory[3837] = 6'd31;
    assign memory[3838] = 6'd32;
    assign memory[3839] = 6'd32;
    assign memory[3840] = 6'd31;
    assign memory[3841] = 6'd31;
    assign memory[3842] = 6'd31;
    assign memory[3843] = 6'd32;
    assign memory[3844] = 6'd32;
    assign memory[3845] = 6'd32;
    assign memory[3846] = 6'd32;
    assign memory[3847] = 6'd31;
    assign memory[3848] = 6'd31;
    assign memory[3849] = 6'd31;
    assign memory[3850] = 6'd32;
    assign memory[3851] = 6'd32;
    assign memory[3852] = 6'd32;
    assign memory[3853] = 6'd32;
    assign memory[3854] = 6'd32;
    assign memory[3855] = 6'd32;
    assign memory[3856] = 6'd32;
    assign memory[3857] = 6'd32;
    assign memory[3858] = 6'd32;
    assign memory[3859] = 6'd31;
    assign memory[3860] = 6'd32;
    assign memory[3861] = 6'd32;
    assign memory[3862] = 6'd32;
    assign memory[3863] = 6'd32;
    assign memory[3864] = 6'd31;
    assign memory[3865] = 6'd31;
    assign memory[3866] = 6'd31;
    assign memory[3867] = 6'd32;
    assign memory[3868] = 6'd32;
    assign memory[3869] = 6'd32;
    assign memory[3870] = 6'd32;
    assign memory[3871] = 6'd32;
    assign memory[3872] = 6'd32;
    assign memory[3873] = 6'd32;
    assign memory[3874] = 6'd31;
    assign memory[3875] = 6'd32;
    assign memory[3876] = 6'd32;
    assign memory[3877] = 6'd32;
    assign memory[3878] = 6'd32;
    assign memory[3879] = 6'd31;
    assign memory[3880] = 6'd32;
    assign memory[3881] = 6'd31;
    assign memory[3882] = 6'd32;
    assign memory[3883] = 6'd32;
    assign memory[3884] = 6'd32;
    assign memory[3885] = 6'd31;
    assign memory[3886] = 6'd31;
    assign memory[3887] = 6'd31;
    assign memory[3888] = 6'd31;
    assign memory[3889] = 6'd32;
    assign memory[3890] = 6'd32;
    assign memory[3891] = 6'd32;
    assign memory[3892] = 6'd32;
    assign memory[3893] = 6'd32;
    assign memory[3894] = 6'd32;
    assign memory[3895] = 6'd31;
    assign memory[3896] = 6'd32;
    assign memory[3897] = 6'd32;
    assign memory[3898] = 6'd31;
    assign memory[3899] = 6'd32;
    assign memory[3900] = 6'd32;
    assign memory[3901] = 6'd32;
    assign memory[3902] = 6'd32;
    assign memory[3903] = 6'd32;
    assign memory[3904] = 6'd32;
    assign memory[3905] = 6'd32;
    assign memory[3906] = 6'd31;
    assign memory[3907] = 6'd32;
    assign memory[3908] = 6'd32;
    assign memory[3909] = 6'd32;
    assign memory[3910] = 6'd32;
    assign memory[3911] = 6'd32;
    assign memory[3912] = 6'd32;
    assign memory[3913] = 6'd32;
    assign memory[3914] = 6'd32;
    assign memory[3915] = 6'd32;
    assign memory[3916] = 6'd31;
    assign memory[3917] = 6'd32;
    assign memory[3918] = 6'd32;
    assign memory[3919] = 6'd32;
    assign memory[3920] = 6'd31;
    assign memory[3921] = 6'd31;
    assign memory[3922] = 6'd32;
    assign memory[3923] = 6'd32;
    assign memory[3924] = 6'd32;
    assign memory[3925] = 6'd32;
    assign memory[3926] = 6'd31;
    assign memory[3927] = 6'd31;
    assign memory[3928] = 6'd31;
    assign memory[3929] = 6'd32;
    assign memory[3930] = 6'd32;
    assign memory[3931] = 6'd32;
    assign memory[3932] = 6'd32;
    assign memory[3933] = 6'd32;
    assign memory[3934] = 6'd32;
    assign memory[3935] = 6'd32;
    assign memory[3936] = 6'd31;
    assign memory[3937] = 6'd32;
    assign memory[3938] = 6'd32;
    assign memory[3939] = 6'd32;
    assign memory[3940] = 6'd32;
    assign memory[3941] = 6'd32;
    assign memory[3942] = 6'd32;
    assign memory[3943] = 6'd31;
    assign memory[3944] = 6'd32;
    assign memory[3945] = 6'd32;
    assign memory[3946] = 6'd32;
    assign memory[3947] = 6'd32;
    assign memory[3948] = 6'd32;
    assign memory[3949] = 6'd32;
    assign memory[3950] = 6'd32;
    assign memory[3951] = 6'd31;
    assign memory[3952] = 6'd31;
    assign memory[3953] = 6'd31;
    assign memory[3954] = 6'd32;
    assign memory[3955] = 6'd33;
    assign memory[3956] = 6'd32;
    assign memory[3957] = 6'd32;
    assign memory[3958] = 6'd32;
    assign memory[3959] = 6'd32;
    assign memory[3960] = 6'd32;
    assign memory[3961] = 6'd31;
    assign memory[3962] = 6'd31;
    assign memory[3963] = 6'd31;
    assign memory[3964] = 6'd32;
    assign memory[3965] = 6'd32;
    assign memory[3966] = 6'd32;
    assign memory[3967] = 6'd31;
    assign memory[3968] = 6'd32;
    assign memory[3969] = 6'd32;
    assign memory[3970] = 6'd32;
    assign memory[3971] = 6'd32;
    assign memory[3972] = 6'd32;
    assign memory[3973] = 6'd31;
    assign memory[3974] = 6'd31;
    assign memory[3975] = 6'd32;
    assign memory[3976] = 6'd31;
    assign memory[3977] = 6'd32;
    assign memory[3978] = 6'd31;
    assign memory[3979] = 6'd32;
    assign memory[3980] = 6'd32;
    assign memory[3981] = 6'd32;
    assign memory[3982] = 6'd32;
    assign memory[3983] = 6'd32;
    assign memory[3984] = 6'd32;
    assign memory[3985] = 6'd31;
    assign memory[3986] = 6'd31;
    assign memory[3987] = 6'd32;
    assign memory[3988] = 6'd32;
    assign memory[3989] = 6'd32;
    assign memory[3990] = 6'd32;
    assign memory[3991] = 6'd32;
    assign memory[3992] = 6'd32;
    assign memory[3993] = 6'd31;
    assign memory[3994] = 6'd32;
    assign memory[3995] = 6'd31;
    assign memory[3996] = 6'd32;
    assign memory[3997] = 6'd31;
    assign memory[3998] = 6'd32;
    assign memory[3999] = 6'd31;
    assign memory[4000] = 6'd31;
    assign memory[4001] = 6'd31;
    assign memory[4002] = 6'd32;
    assign memory[4003] = 6'd32;
    assign memory[4004] = 6'd31;
    assign memory[4005] = 6'd32;
    assign memory[4006] = 6'd31;
    assign memory[4007] = 6'd32;
    assign memory[4008] = 6'd31;
    assign memory[4009] = 6'd32;
    assign memory[4010] = 6'd31;
    assign memory[4011] = 6'd32;
    assign memory[4012] = 6'd32;
    assign memory[4013] = 6'd32;
    assign memory[4014] = 6'd31;
    assign memory[4015] = 6'd32;
    assign memory[4016] = 6'd32;
    assign memory[4017] = 6'd31;
    assign memory[4018] = 6'd32;
    assign memory[4019] = 6'd32;
    assign memory[4020] = 6'd31;
    assign memory[4021] = 6'd32;
    assign memory[4022] = 6'd32;
    assign memory[4023] = 6'd32;
    assign memory[4024] = 6'd32;
    assign memory[4025] = 6'd32;
    assign memory[4026] = 6'd32;
    assign memory[4027] = 6'd32;
    assign memory[4028] = 6'd32;
    assign memory[4029] = 6'd32;
    assign memory[4030] = 6'd32;
    assign memory[4031] = 6'd32;
    assign memory[4032] = 6'd32;
    assign memory[4033] = 6'd31;
    assign memory[4034] = 6'd32;
    assign memory[4035] = 6'd31;
    assign memory[4036] = 6'd32;
    assign memory[4037] = 6'd32;
    assign memory[4038] = 6'd32;
    assign memory[4039] = 6'd32;
    assign memory[4040] = 6'd32;
    assign memory[4041] = 6'd32;
    assign memory[4042] = 6'd32;
    assign memory[4043] = 6'd32;
    assign memory[4044] = 6'd32;
    assign memory[4045] = 6'd32;
    assign memory[4046] = 6'd32;
    assign memory[4047] = 6'd32;
    assign memory[4048] = 6'd32;
    assign memory[4049] = 6'd31;
    assign memory[4050] = 6'd32;
    assign memory[4051] = 6'd31;
    assign memory[4052] = 6'd32;
    assign memory[4053] = 6'd32;
    assign memory[4054] = 6'd32;
    assign memory[4055] = 6'd32;
    assign memory[4056] = 6'd31;
    assign memory[4057] = 6'd32;
    assign memory[4058] = 6'd32;
    assign memory[4059] = 6'd32;
    assign memory[4060] = 6'd32;
    assign memory[4061] = 6'd31;
    assign memory[4062] = 6'd31;
    assign memory[4063] = 6'd32;
    assign memory[4064] = 6'd32;
    assign memory[4065] = 6'd32;
    assign memory[4066] = 6'd32;
    assign memory[4067] = 6'd32;
    assign memory[4068] = 6'd32;
    assign memory[4069] = 6'd32;
    assign memory[4070] = 6'd31;
    assign memory[4071] = 6'd32;
    assign memory[4072] = 6'd31;
    assign memory[4073] = 6'd32;
    assign memory[4074] = 6'd32;
    assign memory[4075] = 6'd31;
    assign memory[4076] = 6'd32;
    assign memory[4077] = 6'd32;
    assign memory[4078] = 6'd32;
    assign memory[4079] = 6'd32;
    assign memory[4080] = 6'd32;
    assign memory[4081] = 6'd32;
    assign memory[4082] = 6'd32;
    assign memory[4083] = 6'd31;
    assign memory[4084] = 6'd31;
    assign memory[4085] = 6'd31;
    assign memory[4086] = 6'd31;
    assign memory[4087] = 6'd32;
    assign memory[4088] = 6'd32;
    assign memory[4089] = 6'd32;
    assign memory[4090] = 6'd32;
    assign memory[4091] = 6'd32;
    assign memory[4092] = 6'd32;
    assign memory[4093] = 6'd32;
    assign memory[4094] = 6'd32;
    assign memory[4095] = 6'd31;

endmodule
