//	How to use:	
//	1. Edit the songs on the Enter Song sheet.	
// 	2. Select this whole worksheet, copy it, and paste it into a new file.	
//	3. Save the file as song_rom.v.	

module pulse5_rom (
    input clk,						
	output reg [25:0] dout,						
	input [11:0] addr		
    );
        
    wire [25:0] memory [4095:0];  				
	always @(posedge clk)						
		dout = memory[addr];					

    parameter s1 = 656;
    parameter s2 = s1 + 120;
    parameter s3 = s2 + 125;

    assign memory[0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[43 ] = {7'd0  , 8'd138, 7'd0  , 2'd0, 2'd0};
    assign memory[44 ] = {7'd30 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4D
    assign memory[45 ] = {7'd33 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4F
    assign memory[46 ] = {7'd35 , 8'd9  , 7'd100, 2'd3, 2'd0};   //note: 4G
    assign memory[47 ] = {7'd37 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4A
    assign memory[48 ] = {7'd38 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[49 ] = {7'd40 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5C
    assign memory[50 ] = {7'd42 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5D
    assign memory[51 ] = {7'd45 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5F
    assign memory[52 ] = {7'd47 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5G
    assign memory[53 ] = {7'd49 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5A
    assign memory[54 ] = {7'd50 , 8'd9  , 7'd100, 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[55 ] = {7'd52 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 6C
    assign memory[56 ] = {7'd54 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[57 ] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[58 ] = {7'd66 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 7D
    assign memory[59 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[60 ] = {7'd59 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[61 ] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[62 ] = {7'd52 , 8'd11 , 7'd96 , 2'd3, 2'd0};   //note: 6C
    assign memory[63 ] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[64 ] = {7'd59 , 8'd11 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[65 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[66 ] = {7'd64 , 8'd13 , 7'd96 , 2'd3, 2'd0};   //note: 7C
    assign memory[67 ] = {7'd0  , 8'd11 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[68 ] = {7'd57 , 8'd13 , 7'd96 , 2'd3, 2'd0};   //note: 6F
    assign memory[69 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[70 ] = {7'd50 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[71 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[72 ] = {7'd57 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 6F
    assign memory[73 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[74 ] = {7'd64 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 7C
    assign memory[75 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[76 ] = {7'd57 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 6F
    assign memory[77 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[78 ] = {7'd50 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[79 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[80 ] = {7'd57 , 8'd13 , 7'd94 , 2'd3, 2'd0};   //note: 6F
    assign memory[81 ] = {7'd0  , 8'd11 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[82 ] = {7'd59 , 8'd13 , 7'd94 , 2'd3, 2'd0};   //note: 6G
    assign memory[83 ] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[84 ] = {7'd55 , 8'd11 , 7'd94 , 2'd3, 2'd0};   //note: 6D#Eb
    assign memory[85 ] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[86 ] = {7'd62 , 8'd11 , 7'd95 , 2'd3, 2'd0};   //note: 6A#Bb
    assign memory[87 ] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[88 ] = {7'd59 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[89 ] = {7'd0  , 8'd10 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[90 ] = {7'd59 , 8'd4  , 7'd121, 2'd3, 2'd0};   //note: 6G
    assign memory[91 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[92 ] = {7'd59 , 8'd4  , 7'd111, 2'd3, 2'd0};   //note: 6G
    assign memory[93 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[94 ] = {7'd59 , 8'd4  , 7'd97 , 2'd3, 2'd0};   //note: 6G
    assign memory[95 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[96 ] = {7'd59 , 8'd4  , 7'd74 , 2'd3, 2'd0};   //note: 6G
    assign memory[97 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[98 ] = {7'd59 , 8'd4  , 7'd57 , 2'd3, 2'd0};   //note: 6G
    assign memory[99 ] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[100] = {7'd59 , 8'd4  , 7'd48 , 2'd3, 2'd0};   //note: 6G
    assign memory[101] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[102] = {7'd59 , 8'd4  , 7'd25 , 2'd3, 2'd0};   //note: 6G
    assign memory[103] = {7'd0  , 8'd44 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[104] = {7'd30 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4D
    assign memory[105] = {7'd33 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4F
    assign memory[106] = {7'd35 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4G
    assign memory[107] = {7'd37 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4A
    assign memory[108] = {7'd40 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5C
    assign memory[109] = {7'd42 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5D
    assign memory[110] = {7'd45 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5F
    assign memory[111] = {7'd47 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5G
    assign memory[112] = {7'd49 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5A
    assign memory[113] = {7'd52 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6C
    assign memory[114] = {7'd54 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[115] = {7'd57 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6F
    assign memory[116] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[117] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[118] = {7'd0  , 8'd162, 7'd0  , 2'd0, 2'd0};
    assign memory[119] = {7'd30 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4D
    assign memory[120] = {7'd33 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4F
    assign memory[121] = {7'd35 , 8'd9  , 7'd100, 2'd3, 2'd0};   //note: 4G
    assign memory[122] = {7'd37 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4A
    assign memory[123] = {7'd38 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[124] = {7'd40 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5C
    assign memory[125] = {7'd42 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5D
    assign memory[126] = {7'd45 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5F
    assign memory[127] = {7'd47 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5G
    assign memory[128] = {7'd49 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5A
    assign memory[129] = {7'd50 , 8'd9  , 7'd100, 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[130] = {7'd52 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 6C
    assign memory[131] = {7'd54 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[132] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[133] = {7'd66 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 7D
    assign memory[134] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[135] = {7'd59 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[136] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[137] = {7'd52 , 8'd11 , 7'd96 , 2'd3, 2'd0};   //note: 6C
    assign memory[138] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[139] = {7'd59 , 8'd11 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[140] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[141] = {7'd64 , 8'd13 , 7'd96 , 2'd3, 2'd0};   //note: 7C
    assign memory[142] = {7'd0  , 8'd11 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[143] = {7'd57 , 8'd13 , 7'd96 , 2'd3, 2'd0};   //note: 6F
    assign memory[144] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[145] = {7'd50 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[146] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[147] = {7'd57 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 6F
    assign memory[148] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[149] = {7'd64 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 7C
    assign memory[150] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[151] = {7'd57 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 6F
    assign memory[152] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[153] = {7'd50 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[154] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[155] = {7'd57 , 8'd13 , 7'd94 , 2'd3, 2'd0};   //note: 6F
    assign memory[156] = {7'd0  , 8'd11 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[157] = {7'd59 , 8'd13 , 7'd94 , 2'd3, 2'd0};   //note: 6G
    assign memory[158] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[159] = {7'd55 , 8'd11 , 7'd94 , 2'd3, 2'd0};   //note: 6D#Eb
    assign memory[160] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[161] = {7'd62 , 8'd11 , 7'd95 , 2'd3, 2'd0};   //note: 6A#Bb
    assign memory[162] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[163] = {7'd59 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[164] = {7'd0  , 8'd10 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[165] = {7'd59 , 8'd4  , 7'd121, 2'd3, 2'd0};   //note: 6G
    assign memory[166] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[167] = {7'd59 , 8'd4  , 7'd111, 2'd3, 2'd0};   //note: 6G
    assign memory[168] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[169] = {7'd59 , 8'd4  , 7'd97 , 2'd3, 2'd0};   //note: 6G
    assign memory[170] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[171] = {7'd59 , 8'd4  , 7'd74 , 2'd3, 2'd0};   //note: 6G
    assign memory[172] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[173] = {7'd59 , 8'd4  , 7'd57 , 2'd3, 2'd0};   //note: 6G
    assign memory[174] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[175] = {7'd59 , 8'd4  , 7'd48 , 2'd3, 2'd0};   //note: 6G
    assign memory[176] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[177] = {7'd59 , 8'd4  , 7'd25 , 2'd3, 2'd0};   //note: 6G
    assign memory[178] = {7'd0  , 8'd44 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[179] = {7'd30 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4D
    assign memory[180] = {7'd33 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4F
    assign memory[181] = {7'd35 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4G
    assign memory[182] = {7'd37 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4A
    assign memory[183] = {7'd40 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5C
    assign memory[184] = {7'd42 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5D
    assign memory[185] = {7'd45 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5F
    assign memory[186] = {7'd47 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5G
    assign memory[187] = {7'd49 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5A
    assign memory[188] = {7'd52 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6C
    assign memory[189] = {7'd54 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[190] = {7'd57 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6F
    assign memory[191] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[192] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[193] = {7'd0  , 8'd162, 7'd0  , 2'd0, 2'd0};
    assign memory[194] = {7'd30 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4D
    assign memory[195] = {7'd33 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4F
    assign memory[196] = {7'd35 , 8'd9  , 7'd100, 2'd3, 2'd0};   //note: 4G
    assign memory[197] = {7'd37 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4A
    assign memory[198] = {7'd38 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[199] = {7'd40 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5C
    assign memory[200] = {7'd42 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5D
    assign memory[201] = {7'd45 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5F
    assign memory[202] = {7'd47 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5G
    assign memory[203] = {7'd49 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5A
    assign memory[204] = {7'd50 , 8'd9  , 7'd100, 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[205] = {7'd52 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 6C
    assign memory[206] = {7'd54 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[207] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[208] = {7'd66 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 7D
    assign memory[209] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[210] = {7'd59 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[211] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[212] = {7'd52 , 8'd11 , 7'd96 , 2'd3, 2'd0};   //note: 6C
    assign memory[213] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[214] = {7'd59 , 8'd11 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[215] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[216] = {7'd64 , 8'd13 , 7'd96 , 2'd3, 2'd0};   //note: 7C
    assign memory[217] = {7'd0  , 8'd11 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[218] = {7'd57 , 8'd13 , 7'd96 , 2'd3, 2'd0};   //note: 6F
    assign memory[219] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[220] = {7'd50 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[221] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[222] = {7'd57 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 6F
    assign memory[223] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[224] = {7'd64 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 7C
    assign memory[225] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[226] = {7'd57 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 6F
    assign memory[227] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[228] = {7'd50 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[229] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[230] = {7'd57 , 8'd13 , 7'd94 , 2'd3, 2'd0};   //note: 6F
    assign memory[231] = {7'd0  , 8'd11 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[232] = {7'd59 , 8'd13 , 7'd94 , 2'd3, 2'd0};   //note: 6G
    assign memory[233] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[234] = {7'd55 , 8'd11 , 7'd94 , 2'd3, 2'd0};   //note: 6D#Eb
    assign memory[235] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[236] = {7'd62 , 8'd11 , 7'd95 , 2'd3, 2'd0};   //note: 6A#Bb
    assign memory[237] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[238] = {7'd59 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[239] = {7'd0  , 8'd10 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[240] = {7'd59 , 8'd4  , 7'd121, 2'd3, 2'd0};   //note: 6G
    assign memory[241] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[242] = {7'd59 , 8'd4  , 7'd111, 2'd3, 2'd0};   //note: 6G
    assign memory[243] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[244] = {7'd59 , 8'd4  , 7'd97 , 2'd3, 2'd0};   //note: 6G
    assign memory[245] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[246] = {7'd59 , 8'd4  , 7'd74 , 2'd3, 2'd0};   //note: 6G
    assign memory[247] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[248] = {7'd59 , 8'd4  , 7'd57 , 2'd3, 2'd0};   //note: 6G
    assign memory[249] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[250] = {7'd59 , 8'd4  , 7'd48 , 2'd3, 2'd0};   //note: 6G
    assign memory[251] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[252] = {7'd59 , 8'd4  , 7'd25 , 2'd3, 2'd0};   //note: 6G
    assign memory[253] = {7'd0  , 8'd44 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[254] = {7'd30 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4D
    assign memory[255] = {7'd33 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4F
    assign memory[256] = {7'd35 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4G
    assign memory[257] = {7'd37 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4A
    assign memory[258] = {7'd40 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5C
    assign memory[259] = {7'd42 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5D
    assign memory[260] = {7'd45 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5F
    assign memory[261] = {7'd47 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5G
    assign memory[262] = {7'd49 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5A
    assign memory[263] = {7'd52 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6C
    assign memory[264] = {7'd54 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[265] = {7'd57 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6F
    assign memory[266] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[267] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[268] = {7'd0  , 8'd162, 7'd0  , 2'd0, 2'd0};
    assign memory[269] = {7'd30 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4D
    assign memory[270] = {7'd33 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4F
    assign memory[271] = {7'd35 , 8'd9  , 7'd100, 2'd3, 2'd0};   //note: 4G
    assign memory[272] = {7'd37 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4A
    assign memory[273] = {7'd38 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[274] = {7'd40 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5C
    assign memory[275] = {7'd42 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5D
    assign memory[276] = {7'd45 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5F
    assign memory[277] = {7'd47 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5G
    assign memory[278] = {7'd49 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 5A
    assign memory[279] = {7'd50 , 8'd9  , 7'd100, 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[280] = {7'd52 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 6C
    assign memory[281] = {7'd54 , 8'd7  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[282] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[283] = {7'd66 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 7D
    assign memory[284] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[285] = {7'd59 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[286] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[287] = {7'd52 , 8'd11 , 7'd96 , 2'd3, 2'd0};   //note: 6C
    assign memory[288] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[289] = {7'd59 , 8'd11 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[290] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[291] = {7'd64 , 8'd13 , 7'd96 , 2'd3, 2'd0};   //note: 7C
    assign memory[292] = {7'd0  , 8'd11 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[293] = {7'd57 , 8'd13 , 7'd96 , 2'd3, 2'd0};   //note: 6F
    assign memory[294] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[295] = {7'd50 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[296] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[297] = {7'd57 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 6F
    assign memory[298] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[299] = {7'd64 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 7C
    assign memory[300] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[301] = {7'd57 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 6F
    assign memory[302] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[303] = {7'd50 , 8'd12 , 7'd95 , 2'd3, 2'd0};   //note: 5A#Bb
    assign memory[304] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[305] = {7'd57 , 8'd13 , 7'd94 , 2'd3, 2'd0};   //note: 6F
    assign memory[306] = {7'd0  , 8'd11 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[307] = {7'd59 , 8'd13 , 7'd94 , 2'd3, 2'd0};   //note: 6G
    assign memory[308] = {7'd0  , 8'd12 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[309] = {7'd55 , 8'd11 , 7'd94 , 2'd3, 2'd0};   //note: 6D#Eb
    assign memory[310] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[311] = {7'd62 , 8'd11 , 7'd95 , 2'd3, 2'd0};   //note: 6A#Bb
    assign memory[312] = {7'd0  , 8'd13 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[313] = {7'd59 , 8'd12 , 7'd96 , 2'd3, 2'd0};   //note: 6G
    assign memory[314] = {7'd0  , 8'd10 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[315] = {7'd59 , 8'd4  , 7'd121, 2'd3, 2'd0};   //note: 6G
    assign memory[316] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[317] = {7'd59 , 8'd4  , 7'd111, 2'd3, 2'd0};   //note: 6G
    assign memory[318] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[319] = {7'd59 , 8'd4  , 7'd97 , 2'd3, 2'd0};   //note: 6G
    assign memory[320] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[321] = {7'd59 , 8'd4  , 7'd74 , 2'd3, 2'd0};   //note: 6G
    assign memory[322] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[323] = {7'd59 , 8'd4  , 7'd57 , 2'd3, 2'd0};   //note: 6G
    assign memory[324] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[325] = {7'd59 , 8'd4  , 7'd48 , 2'd3, 2'd0};   //note: 6G
    assign memory[326] = {7'd0  , 8'd4  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[327] = {7'd59 , 8'd4  , 7'd25 , 2'd3, 2'd0};   //note: 6G
    assign memory[328] = {7'd0  , 8'd44 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[329] = {7'd30 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4D
    assign memory[330] = {7'd33 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4F
    assign memory[331] = {7'd35 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4G
    assign memory[332] = {7'd37 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 4A
    assign memory[333] = {7'd40 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5C
    assign memory[334] = {7'd42 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5D
    assign memory[335] = {7'd45 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5F
    assign memory[336] = {7'd47 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5G
    assign memory[337] = {7'd49 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 5A
    assign memory[338] = {7'd52 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6C
    assign memory[339] = {7'd54 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6D
    assign memory[340] = {7'd57 , 8'd8  , 7'd100, 2'd3, 2'd0};   //note: 6F
    assign memory[341] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[342] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[343] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[344] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[345] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[346] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[347] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[348] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[349] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[350] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[351] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[352] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[353] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[354] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[355] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[356] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[357] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[358] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[359] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[360] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[361] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[362] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[363] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[364] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[365] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[366] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[367] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[368] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[369] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[370] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[371] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[372] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[373] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[374] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[375] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[376] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[377] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[378] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[379] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[380] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[381] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[382] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[383] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[384] = {7'd0  , 8'd171, 7'd0  , 2'd0, 2'd0};
    assign memory[385] = {7'd32 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4E
    assign memory[386] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[387] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[388] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[389] = {7'd32 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4E
    assign memory[390] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[391] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[392] = {7'd0  , 8'd24 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[393] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[394] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[395] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[396] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[397] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[398] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[399] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[400] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[401] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[402] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[403] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[404] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[405] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[406] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[407] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[408] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[409] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[410] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[411] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[412] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[413] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[414] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[415] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[416] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[417] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[418] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[419] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[420] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[421] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[422] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[423] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[424] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[425] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[426] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[427] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[428] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[429] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[430] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[431] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[432] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[433] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[434] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[435] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[436] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[437] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[438] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[439] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[440] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[441] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[442] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[443] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[444] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[445] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[446] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[447] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[448] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[449] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[450] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[451] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[452] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[453] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[454] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[455] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[456] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[457] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[458] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[459] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[460] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[461] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[462] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[463] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[464] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[465] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[466] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[467] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[468] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[469] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[470] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[471] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[472] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[473] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[474] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[475] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[476] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[477] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[478] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[479] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[480] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[481] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[482] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[483] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[484] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[485] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[486] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[487] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[488] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[489] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[490] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[491] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[492] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[493] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[494] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[495] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[496] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[497] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[498] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[499] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[500] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[501] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[502] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[503] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[504] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[505] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[506] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[507] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[508] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[509] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[510] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[511] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[512] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[513] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[514] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[515] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[516] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[517] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[518] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[519] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[520] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[521] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[522] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[523] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[524] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[525] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[526] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[527] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[528] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[529] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[530] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[531] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[532] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[533] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[534] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[535] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[536] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[537] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[538] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[539] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[540] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[541] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[542] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[543] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[544] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[545] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[546] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[547] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[548] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[549] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[550] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[551] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[552] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[553] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[554] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[555] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[556] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[557] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[558] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[559] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[560] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[561] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[562] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[563] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[564] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[565] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[566] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[567] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[568] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[569] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[570] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[571] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[572] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[573] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[574] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[575] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[576] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[577] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[578] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[579] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[580] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[581] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[582] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[583] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[584] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[585] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[586] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[587] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[588] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[589] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[590] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[591] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[592] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[593] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[594] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[595] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[596] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[597] = {7'd33 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4F
    assign memory[598] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[599] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[600] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[601] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[602] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[603] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[604] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[605] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[606] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[607] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[608] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[609] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[610] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[611] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[612] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[613] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[614] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[615] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[616] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[617] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[618] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[619] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[620] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[621] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[622] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[623] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[624] = {7'd45 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5F
    assign memory[625] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[626] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[627] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[628] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[629] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[630] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[631] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[632] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[633] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[634] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[635] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[636] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[637] = {7'd35 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4G
    assign memory[638] = {7'd38 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A#Bb
    assign memory[639] = {7'd42 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5D
    assign memory[640] = {7'd47 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5G
    assign memory[641] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[642] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[643] = {7'd44 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5E
    assign memory[644] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[645] = {7'd37 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 4A
    assign memory[646] = {7'd40 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5C
    assign memory[647] = {7'd44 , 8'd24 , 7'd126, 2'd3, 2'd0};   //note: 5E
    assign memory[648] = {7'd49 , 8'd24 , 7'd127, 2'd3, 2'd0};   //note: 5A
    assign memory[649] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[650] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[651] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[652] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[653] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[654] = {7'd0  , 8'd117, 7'd0  , 2'd0, 2'd0};
    assign memory[655] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s1+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s1+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s1+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+7  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+8  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+9  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+10 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+12 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+13 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+14 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+15 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+16 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+17 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+18 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+19 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+20 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+21 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+22 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+23 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+24 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+25 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+26 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+27 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+28 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+29 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+30 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+31 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+32 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+33 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+34 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+35 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+36 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+37 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+38 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+45 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+46 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+47 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+48 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+49 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+50 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+51 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+52 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+53 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+54 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+55 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+56 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+57 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+58 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+59 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+60 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+61 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+62 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+63 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+64 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+65 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+66 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+67 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+68 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+69 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+70 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+71 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+72 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+73 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+74 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+75 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+76 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+77 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+78 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+79 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+80 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+81 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+82 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+83 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+84 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+85 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+86 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+87 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+88 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+89 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+90 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+91 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+92 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+93 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+94 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+95 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+96 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+97 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+98 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+99 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+100] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+101] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+102] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+103] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+104] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+105] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+106] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+107] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+108] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+109] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+110] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+111] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+112] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+113] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+114] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+115] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+116] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+117] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+118] = {7'd0  , 8'd118, 7'd0  , 2'd0, 2'd0};
    assign memory[s1+119] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s2+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s2+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+2  ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+3  ] = {7'd33 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+4  ] = {7'd33 , 8'd129, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+5  ] = {7'd29 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+6  ] = {7'd29 , 8'd129, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+7  ] = {7'd31 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+8  ] = {7'd31 , 8'd129, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+9  ] = {7'd31 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+10 ] = {7'd31 , 8'd129, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+11 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+12 ] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+13 ] = {7'd28 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4C
    assign memory[s2+14 ] = {7'd28 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+15 ] = {7'd29 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+16 ] = {7'd29 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+17 ] = {7'd24 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 3G#Ab
    assign memory[s2+18 ] = {7'd24 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+19 ] = {7'd26 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s2+20 ] = {7'd26 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+21 ] = {7'd28 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4C
    assign memory[s2+22 ] = {7'd28 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+23 ] = {7'd29 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+24 ] = {7'd29 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+25 ] = {7'd24 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 3G#Ab
    assign memory[s2+26 ] = {7'd24 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+27 ] = {7'd26 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 3A#Bb
    assign memory[s2+28 ] = {7'd26 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+29 ] = {7'd33 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+30 ] = {7'd33 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+31 ] = {7'd29 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+32 ] = {7'd29 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+33 ] = {7'd31 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+34 ] = {7'd31 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+35 ] = {7'd31 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+36 ] = {7'd31 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+37 ] = {7'd33 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+38 ] = {7'd33 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+39 ] = {7'd29 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+40 ] = {7'd29 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+41 ] = {7'd31 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+42 ] = {7'd31 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+43 ] = {7'd31 , 8'd255, 7'd80 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+44 ] = {7'd31 , 8'd129, 7'd80 , 2'd0, 2'd0};
    assign memory[s2+45 ] = {7'd33 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+46 ] = {7'd33 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+47 ] = {7'd36 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+48 ] = {7'd36 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+49 ] = {7'd31 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+50 ] = {7'd31 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+51 ] = {7'd35 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 4G
    assign memory[s2+52 ] = {7'd35 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+53 ] = {7'd33 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+54 ] = {7'd33 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+55 ] = {7'd36 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+56 ] = {7'd36 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+57 ] = {7'd36 , 8'd255, 7'd95 , 2'd0, 2'd0};   //note: 4G#Ab
    assign memory[s2+58 ] = {7'd36 , 8'd129, 7'd95 , 2'd0, 2'd0};
    assign memory[s2+59 ] = {7'd35 , 8'd192, 7'd95 , 2'd0, 2'd0};   //note: 4G
    assign memory[s2+60 ] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+61 ] = {7'd33 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4F
    assign memory[s2+62 ] = {7'd33 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+63 ] = {7'd33 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4F
    assign memory[s2+64 ] = {7'd29 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+65 ] = {7'd29 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+66 ] = {7'd29 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+67 ] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+68 ] = {7'd31 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+69 ] = {7'd31 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+70 ] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+71 ] = {7'd31 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+72 ] = {7'd31 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+73 ] = {7'd33 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4F
    assign memory[s2+74 ] = {7'd33 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+75 ] = {7'd33 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4F
    assign memory[s2+76 ] = {7'd29 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+77 ] = {7'd29 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+78 ] = {7'd29 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+79 ] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+80 ] = {7'd31 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+81 ] = {7'd31 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+82 ] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+83 ] = {7'd31 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+84 ] = {7'd31 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+85 ] = {7'd33 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4F
    assign memory[s2+86 ] = {7'd33 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+87 ] = {7'd33 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4F
    assign memory[s2+88 ] = {7'd29 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+89 ] = {7'd29 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+90 ] = {7'd29 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+91 ] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+92 ] = {7'd31 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+93 ] = {7'd31 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+94 ] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+95 ] = {7'd31 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+96 ] = {7'd31 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+97 ] = {7'd33 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4F
    assign memory[s2+98 ] = {7'd33 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+99 ] = {7'd33 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4F
    assign memory[s2+100] = {7'd29 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+101] = {7'd29 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+102] = {7'd29 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+103] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+104] = {7'd31 , 8'd33 , 7'd100, 2'd0, 2'd0};
    assign memory[s2+105] = {7'd31 , 8'd96 , 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+106] = {7'd31 , 8'd255, 7'd100, 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+107] = {7'd31 , 8'd129, 7'd100, 2'd0, 2'd0};
    assign memory[s2+108] = {7'd33 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+109] = {7'd33 , 8'd33 , 7'd72 , 2'd0, 2'd0};
    assign memory[s2+110] = {7'd33 , 8'd96 , 7'd72 , 2'd0, 2'd0};   //note: 4F
    assign memory[s2+111] = {7'd29 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+112] = {7'd29 , 8'd33 , 7'd72 , 2'd0, 2'd0};
    assign memory[s2+113] = {7'd29 , 8'd96 , 7'd72 , 2'd0, 2'd0};   //note: 4C#Db
    assign memory[s2+114] = {7'd31 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+115] = {7'd31 , 8'd33 , 7'd72 , 2'd0, 2'd0};
    assign memory[s2+116] = {7'd31 , 8'd96 , 7'd72 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+117] = {7'd31 , 8'd255, 7'd72 , 2'd0, 2'd0};   //note: 4D#Eb
    assign memory[s2+118] = {7'd31 , 8'd255, 7'd72 , 2'd0, 2'd0};
    assign memory[s2+119] = {7'd31 , 8'd66 , 7'd72 , 2'd0, 2'd0};
    assign memory[s2+120] = {7'd0  , 8'd192, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+121] = {7'd0  , 8'd1  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+122] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s2+123] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s2+124] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song

    assign memory[s3+0  ] = {7'd126, 8'd0  , 7'd0  , 2'd0, 2'd0};   //Begin of a song
    assign memory[s3+1  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+2  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+3  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+4  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+5  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+6  ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+7  ] = {7'd0  , 8'd102, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+8  ] = {7'd24 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+9  ] = {7'd27 , 8'd24 , 7'd79 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+10 ] = {7'd31 , 8'd72 , 7'd79 , 2'd2, 2'd0};   //note: 4D#Eb
    assign memory[s3+11 ] = {7'd27 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+12 ] = {7'd22 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+13 ] = {7'd26 , 8'd24 , 7'd79 , 2'd2, 2'd0};   //note: 3A#Bb
    assign memory[s3+14 ] = {7'd29 , 8'd72 , 7'd79 , 2'd2, 2'd0};   //note: 4C#Db
    assign memory[s3+15 ] = {7'd26 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3A#Bb
    assign memory[s3+16 ] = {7'd20 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+17 ] = {7'd24 , 8'd24 , 7'd79 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+18 ] = {7'd27 , 8'd72 , 7'd79 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+19 ] = {7'd24 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+20 ] = {7'd15 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+21 ] = {7'd19 , 8'd24 , 7'd79 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+22 ] = {7'd22 , 8'd72 , 7'd79 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+23 ] = {7'd19 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+24 ] = {7'd15 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+25 ] = {7'd20 , 8'd24 , 7'd79 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+26 ] = {7'd22 , 8'd72 , 7'd79 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+27 ] = {7'd20 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+28 ] = {7'd19 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+29 ] = {7'd22 , 8'd24 , 7'd79 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+30 ] = {7'd27 , 8'd72 , 7'd79 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+31 ] = {7'd22 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+32 ] = {7'd22 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+33 ] = {7'd26 , 8'd24 , 7'd79 , 2'd2, 2'd0};   //note: 3A#Bb
    assign memory[s3+34 ] = {7'd29 , 8'd72 , 7'd79 , 2'd2, 2'd0};   //note: 4C#Db
    assign memory[s3+35 ] = {7'd26 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3A#Bb
    assign memory[s3+36 ] = {7'd27 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+37 ] = {7'd22 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+38 ] = {7'd27 , 8'd48 , 7'd79 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+39 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+40 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+41 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+42 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+43 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+44 ] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+45 ] = {7'd0  , 8'd54 , 7'd0  , 2'd0, 2'd0};
    assign memory[s3+46 ] = {7'd20 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+47 ] = {7'd20 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+48 ] = {7'd27 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+49 ] = {7'd20 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+50 ] = {7'd15 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+51 ] = {7'd15 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+52 ] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+53 ] = {7'd15 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+54 ] = {7'd10 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 2F#Gb
    assign memory[s3+55 ] = {7'd10 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 2F#Gb
    assign memory[s3+56 ] = {7'd17 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3C#Db
    assign memory[s3+57 ] = {7'd10 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 2F#Gb
    assign memory[s3+58 ] = {7'd12 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 2G#Ab
    assign memory[s3+59 ] = {7'd12 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 2G#Ab
    assign memory[s3+60 ] = {7'd19 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+61 ] = {7'd12 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 2G#Ab
    assign memory[s3+62 ] = {7'd20 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+63 ] = {7'd20 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+64 ] = {7'd27 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+65 ] = {7'd20 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+66 ] = {7'd15 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+67 ] = {7'd15 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+68 ] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+69 ] = {7'd15 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+70 ] = {7'd22 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+71 ] = {7'd22 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+72 ] = {7'd29 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 4C#Db
    assign memory[s3+73 ] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+74 ] = {7'd23 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+75 ] = {7'd23 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+76 ] = {7'd29 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 4C#Db
    assign memory[s3+77 ] = {7'd23 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+78 ] = {7'd20 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+79 ] = {7'd20 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+80 ] = {7'd27 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+81 ] = {7'd20 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+82 ] = {7'd15 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+83 ] = {7'd15 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+84 ] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+85 ] = {7'd15 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+86 ] = {7'd19 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+87 ] = {7'd19 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+88 ] = {7'd23 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+89 ] = {7'd19 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+90 ] = {7'd24 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+91 ] = {7'd24 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+92 ] = {7'd31 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 4D#Eb
    assign memory[s3+93 ] = {7'd24 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+94 ] = {7'd20 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+95 ] = {7'd20 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+96 ] = {7'd27 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+97 ] = {7'd20 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+98 ] = {7'd19 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+99 ] = {7'd19 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+100] = {7'd27 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+101] = {7'd19 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+102] = {7'd20 , 8'd96 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+103] = {7'd22 , 8'd96 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+104] = {7'd21 , 8'd96 , 7'd99 , 2'd2, 2'd0};   //note: 3F
    assign memory[s3+105] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+106] = {7'd20 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+107] = {7'd20 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+108] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+109] = {7'd20 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+110] = {7'd19 , 8'd72 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+111] = {7'd19 , 8'd24 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+112] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+113] = {7'd19 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+114] = {7'd20 , 8'd96 , 7'd99 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+115] = {7'd22 , 8'd96 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+116] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+117] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+118] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+119] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+120] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+121] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+122] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+123] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+124] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+125] = {7'd22 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+126] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+127] = {7'd23 , 8'd48 , 7'd99 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+128] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+129] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+130] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+131] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+132] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+133] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+134] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+135] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+136] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+137] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+138] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+139] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+140] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+141] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+142] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+143] = {7'd0  , 8'd87 , 7'd0  , 2'd0, 2'd0};
    assign memory[s3+144] = {7'd20 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+145] = {7'd27 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+146] = {7'd20 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+147] = {7'd15 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+148] = {7'd15 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+149] = {7'd22 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+150] = {7'd15 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+151] = {7'd10 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 2F#Gb
    assign memory[s3+152] = {7'd10 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 2F#Gb
    assign memory[s3+153] = {7'd17 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3C#Db
    assign memory[s3+154] = {7'd10 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 2F#Gb
    assign memory[s3+155] = {7'd12 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 2G#Ab
    assign memory[s3+156] = {7'd12 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 2G#Ab
    assign memory[s3+157] = {7'd19 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+158] = {7'd12 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 2G#Ab
    assign memory[s3+159] = {7'd20 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+160] = {7'd20 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+161] = {7'd27 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+162] = {7'd20 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+163] = {7'd15 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+164] = {7'd15 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+165] = {7'd22 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+166] = {7'd15 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+167] = {7'd22 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+168] = {7'd22 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+169] = {7'd29 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 4C#Db
    assign memory[s3+170] = {7'd22 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+171] = {7'd23 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+172] = {7'd23 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+173] = {7'd29 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 4C#Db
    assign memory[s3+174] = {7'd23 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+175] = {7'd20 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+176] = {7'd20 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+177] = {7'd27 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+178] = {7'd20 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+179] = {7'd15 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+180] = {7'd15 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+181] = {7'd22 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+182] = {7'd15 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 2B
    assign memory[s3+183] = {7'd19 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+184] = {7'd19 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+185] = {7'd23 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3G
    assign memory[s3+186] = {7'd19 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+187] = {7'd24 , 8'd72 , 7'd94 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+188] = {7'd24 , 8'd24 , 7'd94 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+189] = {7'd31 , 8'd48 , 7'd94 , 2'd2, 2'd0};   //note: 4D#Eb
    assign memory[s3+190] = {7'd24 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3G#Ab
    assign memory[s3+191] = {7'd20 , 8'd72 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+192] = {7'd20 , 8'd24 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+193] = {7'd27 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+194] = {7'd20 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+195] = {7'd19 , 8'd72 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+196] = {7'd19 , 8'd24 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+197] = {7'd27 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3B
    assign memory[s3+198] = {7'd19 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+199] = {7'd20 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+200] = {7'd22 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+201] = {7'd21 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3F
    assign memory[s3+202] = {7'd0  , 8'd96 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+203] = {7'd20 , 8'd72 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+204] = {7'd20 , 8'd24 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+205] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+206] = {7'd20 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+207] = {7'd19 , 8'd72 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+208] = {7'd19 , 8'd24 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+209] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+210] = {7'd19 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+211] = {7'd20 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+212] = {7'd22 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+213] = {7'd22 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+214] = {7'd19 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+215] = {7'd20 , 8'd72 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+216] = {7'd20 , 8'd24 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+217] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+218] = {7'd20 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+219] = {7'd19 , 8'd72 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+220] = {7'd19 , 8'd24 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+221] = {7'd0  , 8'd48 , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+222] = {7'd19 , 8'd48 , 7'd95 , 2'd2, 2'd0};   //note: 3D#Eb
    assign memory[s3+223] = {7'd20 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3E
    assign memory[s3+224] = {7'd22 , 8'd96 , 7'd95 , 2'd2, 2'd0};   //note: 3F#Gb
    assign memory[s3+225] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+226] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+227] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+228] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+229] = {7'd0  , 8'd132, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+230] = {7'd0  , 8'd2  , 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+231] = {7'd0  , 8'd255, 7'd0  , 2'd0, 2'd0};   //note: rest
    assign memory[s3+232] = {7'd0  , 8'd129, 7'd0  , 2'd0, 2'd0};
    assign memory[s3+233] = {7'd127, 8'd0  , 7'd0  , 2'd0, 2'd0};   //End of a song


endmodule							
